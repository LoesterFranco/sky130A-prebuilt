* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_80_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=6.012e+11p ps=5.38e+06u
M1001 a_356_392# B1 a_80_392# VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1002 a_168_136# A1 a_85_136# VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=5.184e+11p ps=5.46e+06u
M1003 a_85_136# D1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=7.465e+11p ps=6.29e+06u
M1004 a_85_136# D1 a_434_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1005 VGND A2 a_168_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_85_136# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C1 a_85_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_85_136# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1009 a_434_392# C1 a_356_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_80_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_85_136# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_633_368# B1 a_525_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.944e+11p pd=5.72e+06u as=4.032e+11p ps=2.96e+06u
M1001 a_447_368# D1 a_91_244# VPB pshort w=1.12e+06u l=180000u
+  ad=2.352e+11p pd=2.66e+06u as=2.912e+11p ps=2.76e+06u
M1002 VPWR A2 a_633_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.856e+11p pd=8.48e+06u as=0p ps=0u
M1003 a_91_244# C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=1.0508e+12p ps=8.76e+06u
M1004 X a_91_244# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VPWR a_91_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_525_368# C1 a_447_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_633_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_91_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1009 X a_91_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_771_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1011 a_91_244# A1 a_771_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B1 a_91_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D1 a_91_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_1013_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.06e+12p pd=1.012e+07u as=1.4248e+12p ps=1.338e+07u
M1001 a_137_260# A1 a_1210_74# VNB nlowvt w=640000u l=150000u
+  ad=7.168e+11p pd=7.36e+06u as=5.184e+11p ps=5.46e+06u
M1002 a_137_260# D1 a_549_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u
M1003 VGND a_137_260# X VNB nlowvt w=740000u l=150000u
+  ad=1.3711e+12p pd=1.359e+07u as=4.144e+11p ps=4.08e+06u
M1004 VGND C1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_549_392# D1 a_137_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_817_392# C1 a_549_392# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1007 a_1210_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_549_392# C1 a_817_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_137_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_137_260# D1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1210_74# A1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_817_392# B1 a_1013_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_137_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1015 a_1013_392# B1 a_817_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_137_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_1013_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_137_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1013_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_137_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND D1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_137_260# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_137_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_137_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A2 a_1013_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_137_260# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_1210_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_345_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.944e+11p pd=5.72e+06u as=4.032e+11p ps=2.96e+06u
M1001 VGND A2 a_461_74# VNB nlowvt w=740000u l=150000u
+  ad=7.77e+11p pd=6.54e+06u as=2.368e+11p ps=2.12e+06u
M1002 a_461_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1003 Y D1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_237_368# C1 a_159_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=2.352e+11p ps=2.66e+06u
M1005 a_345_368# B1 a_237_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_159_368# D1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1008 VPWR A1 a_345_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=7.141e+11p pd=6.37e+06u as=6.919e+11p ps=6.31e+06u
M1001 a_722_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=0p ps=0u
M1002 a_533_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.1872e+12p pd=1.108e+07u as=6.048e+11p ps=5.56e+06u
M1003 Y D1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=8.848e+11p ps=8.3e+06u
M1004 a_69_368# D1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_722_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_337_368# C1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1007 Y D1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_69_368# C1 a_337_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_337_368# B1 a_533_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_533_368# B1 a_337_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A1 a_533_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_722_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A1 a_722_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_533_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A2 a_533_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_477_368# C1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=1.4896e+12p ps=1.386e+07u
M1001 VPWR A1 a_853_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=2.1168e+12p ps=1.946e+07u
M1002 a_29_368# C1 a_477_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_853_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_477_368# C1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_853_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_29_368# C1 a_477_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_1228_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0434e+12p pd=1.022e+07u as=1.887e+12p ps=1.398e+07u
M1008 a_853_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1228_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.036e+12p ps=1.02e+07u
M1010 VPWR A2 a_853_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1228_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_477_368# B1 a_853_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_853_368# B1 a_477_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_853_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y D1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A2 a_1228_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_477_368# B1 a_853_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y D1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1022 a_29_368# D1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1228_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_853_368# B1 a_477_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y D1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_1228_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR A1 a_853_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND D1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A1 a_1228_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_29_368# D1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_853_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y A1 a_1228_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VGND a_81_264# X VNB nlowvt w=740000u l=150000u
+  ad=5.3685e+11p pd=4.68e+06u as=1.961e+11p ps=2.01e+06u
M1001 a_81_264# C1 a_553_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1002 a_279_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=5.912e+11p ps=5.36e+06u
M1003 VGND B1 a_81_264# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.488e+11p ps=3.65e+06u
M1004 a_81_264# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_553_392# B1 a_279_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_366_136# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=2.08e+11p pd=1.93e+06u as=0p ps=0u
M1007 VPWR a_81_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1008 a_81_264# A1 a_366_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_279_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_317_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=9.424e+11p ps=8.24e+06u
M1001 a_85_270# A1 a_399_74# VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=1.554e+11p ps=1.9e+06u
M1002 a_603_392# B1 a_317_392# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1003 a_399_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=9.731e+11p ps=7.07e+06u
M1004 VGND a_85_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 VGND B1 a_85_270# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_85_270# C1 a_603_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1007 VPWR A2 a_317_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_85_270# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_85_270# C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_85_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1011 VPWR a_85_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_1064_123# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=1.50765e+12p ps=1.284e+07u
M1001 X a_105_280# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1002 a_105_280# A1 a_1064_123# VNB nlowvt w=640000u l=150000u
+  ad=5.79525e+11p pd=5.76e+06u as=0p ps=0u
M1003 VPWR A1 a_517_392# VPB pshort w=1e+06u l=180000u
+  ad=1.7798e+12p pd=1.409e+07u as=1.065e+12p ps=1.013e+07u
M1004 a_517_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_105_280# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_105_280# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1007 VGND a_105_280# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_105_280# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_105_280# C1 a_605_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=6.15e+11p ps=5.23e+06u
M1010 a_605_392# B1 a_517_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_105_280# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_605_392# C1 a_105_280# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B1 a_105_280# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_517_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_105_280# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_105_280# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1064_123# A1 a_105_280# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_517_392# B1 a_605_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_105_280# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_105_280# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND C1 a_105_280# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_517_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A2 a_1064_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_71_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=4.032e+11p ps=2.96e+06u
M1001 Y A1 a_159_74# VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=1.554e+11p ps=1.9e+06u
M1002 a_357_368# B1 a_71_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1003 a_159_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.847e+11p ps=4.27e+06u
M1004 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_71_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 a_357_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1007 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_38_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=6.438e+11p ps=6.18e+06u
M1001 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=7.4e+11p pd=4.96e+06u as=0p ps=0u
M1002 VGND A2 a_38_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_368# B1 a_497_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.072e+11p pd=8.34e+06u as=9.072e+11p ps=8.34e+06u
M1004 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_497_368# B1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 a_497_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1007 Y A1 a_38_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_497_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_38_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_117_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=9.072e+11p ps=8.34e+06u
M1011 VPWR A1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_117_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A2 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_92_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.0286e+12p pd=1.018e+07u as=1.0138e+12p ps=1.014e+07u
M1001 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.288e+11p ps=8.16e+06u
M1002 Y C1 a_901_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.4896e+12p ps=1.386e+07u
M1003 VGND A2 a_92_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_901_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_92_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A2 a_77_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=2.0944e+12p ps=1.942e+07u
M1007 a_77_368# B1 a_901_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A1 a_92_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_77_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_92_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_77_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_92_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_901_368# B1 a_77_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_77_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_77_368# B1 a_901_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A1 a_92_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A1 a_77_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_901_368# B1 a_77_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_77_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y C1 a_901_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_77_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_901_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_77_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_92_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_34_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=6.766e+11p ps=5.55e+06u
M1001 X a_194_136# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1002 a_122_136# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=5.6545e+11p ps=5.75e+06u
M1003 X a_194_136# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1004 VGND a_272_110# a_194_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.496e+11p ps=2.06e+06u
M1005 a_194_136# a_272_110# a_34_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1006 VPWR A2 a_34_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1_N a_272_110# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1008 VGND B1_N a_272_110# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 a_194_136# A1 a_122_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VGND a_187_244# X VNB nlowvt w=740000u l=150000u
+  ad=9.689e+11p pd=7.11e+06u as=2.072e+11p ps=2.04e+06u
M1001 VPWR B1_N a_32_368# VPB pshort w=840000u l=180000u
+  ad=9.154e+11p pd=8.21e+06u as=2.184e+11p ps=2.2e+06u
M1002 X a_187_244# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1003 a_187_244# a_32_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 VPWR a_187_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_187_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_507_392# a_32_368# a_187_244# VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=2.6e+11p ps=2.52e+06u
M1007 VPWR A1 a_507_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_507_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_587_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1010 VGND B1_N a_32_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.4575e+11p ps=1.63e+06u
M1011 a_587_74# A1 a_187_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_184_338# a_29_392# a_596_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.06e+12p ps=1.012e+07u
M1001 VPWR a_184_338# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.4998e+12p pd=1.353e+07u as=6.048e+11p ps=5.56e+06u
M1002 a_596_392# a_29_392# a_184_338# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_184_338# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.34918e+12p ps=1.097e+07u
M1004 X a_184_338# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_596_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_184_338# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_596_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_184_338# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1_N a_29_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1010 a_864_123# A1 a_184_338# VNB nlowvt w=640000u l=150000u
+  ad=3.968e+11p pd=3.8e+06u as=3.584e+11p ps=3.68e+06u
M1011 X a_184_338# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_864_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_184_338# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_184_338# A1 a_864_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_596_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B1_N a_29_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1017 VGND a_29_392# a_184_338# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_596_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_864_123# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_184_338# a_29_392# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_184_338# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_437_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=2.072e+11p ps=2.04e+06u
M1001 VGND B1_N a_29_424# VNB nlowvt w=550000u l=150000u
+  ad=5.5275e+11p pd=4.59e+06u as=1.4575e+11p ps=1.63e+06u
M1002 a_351_368# a_29_424# Y VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=2.912e+11p ps=2.76e+06u
M1003 a_351_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.544e+11p ps=5.04e+06u
M1004 VPWR A1 a_351_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_29_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_437_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1_N a_29_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_436_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=4.144e+11p ps=4.08e+06u
M1001 Y a_62_94# a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1872e+12p ps=1.108e+07u
M1002 a_241_368# a_62_94# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B1_N a_62_94# VNB nlowvt w=640000u l=150000u
+  ad=6.474e+11p pd=6.21e+06u as=1.696e+11p ps=1.81e+06u
M1004 VPWR A1 a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=8.872e+11p pd=8.12e+06u as=0p ps=0u
M1005 a_241_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_62_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_436_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2 a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_241_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_62_94# B1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1011 VGND a_62_94# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A1 a_436_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_436_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VGND a_803_323# Y VNB nlowvt w=740000u l=150000u
+  ad=1.0249e+12p pd=1.017e+07u as=8.288e+11p ps=8.16e+06u
M1001 Y a_803_323# a_31_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=2.0944e+12p ps=1.942e+07u
M1002 a_46_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0138e+12p pd=1.014e+07u as=0p ps=0u
M1003 a_46_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_803_323# B1_N VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1005 Y A1 a_46_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_46_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_31_368# a_803_323# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_31_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.6464e+12p pd=1.552e+07u as=0p ps=0u
M1009 a_31_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_31_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A2 a_46_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_46_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_803_323# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_31_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_46_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A2 a_31_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_803_323# B1_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1018 a_31_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B1_N a_803_323# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A2 a_31_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y a_803_323# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_31_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_46_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_803_323# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y a_803_323# a_31_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_31_368# a_803_323# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VGND a_81_264# X VNB nlowvt w=740000u l=150000u
+  ad=4.541e+11p pd=4.09e+06u as=1.961e+11p ps=2.01e+06u
M1001 VGND A2 a_452_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.93e+06u
M1002 a_367_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=5.912e+11p ps=5.36e+06u
M1003 a_81_264# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1004 a_452_136# A1 a_81_264# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_81_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1006 a_367_392# B1 a_81_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1007 VPWR A1 a_367_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_404_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=8.524e+11p ps=8.06e+06u
M1001 X a_84_244# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1002 VPWR a_84_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_84_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.954e+11p ps=6.86e+06u
M1004 a_84_244# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VGND a_84_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_484_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1007 a_404_392# B1 a_84_244# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1008 a_484_74# A1 a_84_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_404_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_700_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=5.184e+11p pd=5.46e+06u as=1.011e+12p ps=9.9e+06u
M1001 X a_91_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1002 a_503_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.06e+12p pd=1.012e+07u as=1.4248e+12p ps=1.338e+07u
M1003 a_700_74# A1 a_91_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1004 X a_91_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_91_48# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_91_48# B1 a_503_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1007 X a_91_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1008 VPWR a_91_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_503_392# B1 a_91_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_91_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_91_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_91_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_503_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_91_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_700_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_503_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_91_48# A1 a_700_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A2 a_503_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 a_91_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_29_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=3.36e+11p ps=2.84e+06u
M1001 Y B1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1002 Y A1 a_117_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1003 VPWR A2 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.07e+11p pd=4.06e+06u as=0p ps=0u
M1005 a_117_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_280_107# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=6.5505e+11p pd=6.27e+06u as=4.033e+11p ps=4.05e+06u
M1001 a_280_107# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.83425e+11p ps=4.82e+06u
M1002 VGND A2 a_280_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 a_131_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1872e+12p ps=1.108e+07u
M1004 a_131_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_131_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1006 Y A1 a_280_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_131_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_131_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_131_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 Y A1 a_84_74# VNB nlowvt w=740000u l=150000u
+  ad=8.066e+11p pd=8.1e+06u as=1.0286e+12p ps=1.018e+07u
M1001 Y A1 a_84_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_84_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=6.216e+11p ps=6.12e+06u
M1003 VPWR A2 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=2.0944e+12p ps=1.942e+07u
M1004 Y B1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1005 a_69_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_69_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A2 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_69_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_84_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_84_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_69_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_84_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_84_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A2 a_84_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_69_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_69_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VPWR a_148_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=6.262e+11p pd=5.43e+06u as=2.912e+11p ps=2.76e+06u
M1001 a_313_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1002 VPWR A1 a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_148_260# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=4.192e+11p pd=3.87e+06u as=8.64875e+11p ps=5.71e+06u
M1004 a_417_79# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1005 a_148_260# A1 a_417_79# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_148_260# C1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=5.6e+11p ps=5.12e+06u
M1007 VGND a_148_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1008 a_597_79# B1 a_148_260# VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1009 VGND B2 a_597_79# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_313_392# B1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_509_392# B2 a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_319_392# VPB pshort w=1e+06u l=180000u
+  ad=9.174e+11p pd=8.19e+06u as=5.4e+11p ps=5.08e+06u
M1001 a_89_260# A1 a_337_74# VNB nlowvt w=740000u l=150000u
+  ad=8.029e+11p pd=5.13e+06u as=1.554e+11p ps=1.9e+06u
M1002 X a_89_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.362e+11p ps=6.7e+06u
M1003 VGND a_89_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_319_392# B1 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.3e+11p ps=5.06e+06u
M1005 a_515_392# B2 a_319_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_89_260# C1 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1007 a_337_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_603_74# B1 a_89_260# VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1009 VGND B2 a_603_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_89_260# C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_89_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1012 VPWR a_89_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_319_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_1102_392# C1 a_154_135# VPB pshort w=1e+06u l=180000u
+  ad=1.35e+12p pd=1.07e+07u as=2.7e+11p ps=2.54e+06u
M1001 a_160_376# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.24e+12p pd=1.048e+07u as=2.0298e+12p ps=1.459e+07u
M1002 a_160_376# B2 a_1102_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A2 a_160_376# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1102_392# B2 a_160_376# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_154_135# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.62282e+12p ps=1.315e+07u
M1006 X a_154_135# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1007 a_160_376# B1 a_1102_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_154_135# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_154_135# A1 a_71_135# VNB nlowvt w=640000u l=150000u
+  ad=5.376e+11p pd=5.52e+06u as=5.184e+11p ps=5.46e+06u
M1010 X a_154_135# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_71_135# A1 a_154_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_154_135# B1 a_1346_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.632e+11p ps=5.6e+06u
M1013 VPWR a_154_135# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1102_392# B1 a_160_376# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_154_135# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_160_376# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1346_123# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_160_376# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B2 a_1346_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1346_123# B1 a_154_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_154_135# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_71_135# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_154_135# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_154_135# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND C1 a_154_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_154_135# C1 a_1102_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_71_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 Y B1 a_351_74# VNB nlowvt w=740000u l=150000u
+  ad=8.695e+11p pd=5.31e+06u as=1.554e+11p ps=1.9e+06u
M1001 a_121_368# B2 a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=9.184e+11p ps=8.36e+06u
M1002 VPWR A1 a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=0p ps=0u
M1003 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=0p ps=0u
M1004 a_263_368# B1 a_121_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_263_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_567_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1007 VGND A2 a_567_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_351_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_121_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_297_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2432e+12p pd=1.118e+07u as=8.848e+11p ps=8.3e+06u
M1001 VGND B2 a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=7.696e+11p pd=6.52e+06u as=4.44e+11p ps=4.16e+06u
M1002 VPWR A2 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_293_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.362e+11p ps=8.18e+06u
M1004 a_675_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=7.03e+11p pd=4.86e+06u as=0p ps=0u
M1005 a_297_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_675_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_675_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_293_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_29_368# B2 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1872e+12p pd=1.108e+07u as=0p ps=0u
M1011 a_297_368# B2 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_29_368# B1 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_675_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1017 a_29_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_297_368# B1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_117_368# B1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.8144e+12p pd=1.668e+07u as=2.6992e+12p ps=2.498e+07u
M1001 VGND A2 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=1.2432e+12p pd=1.224e+07u as=1.0138e+12p ps=1.014e+07u
M1002 VPWR A2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.4672e+12p pd=1.158e+07u as=0p ps=0u
M1003 a_531_368# B1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1326_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0138e+12p pd=1.014e+07u as=0p ps=0u
M1005 VGND A2 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B2 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_531_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_117_368# B1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1326_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.4282e+12p ps=1.422e+07u
M1010 a_534_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_531_368# B1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1326_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_531_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_117_368# B2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_534_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_531_368# B2 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_534_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1326_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B2 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_117_368# B2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A1 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y B1 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_531_368# B2 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_531_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_117_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=8.848e+11p ps=8.3e+06u
M1032 Y C1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y A1 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_534_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_117_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y B1 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y C1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_531_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a222o_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
M1000 VGND C2 a_119_74# VNB nlowvt w=640000u l=150000u
+  ad=9.082e+11p pd=5.52e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_32_74# C1 a_27_390# VPB pshort w=1e+06u l=180000u
+  ad=4.25e+11p pd=2.85e+06u as=8.8e+11p ps=7.76e+06u
M1002 X a_32_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 VGND A2 a_651_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1004 a_651_74# A1 a_32_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=6.848e+11p ps=4.7e+06u
M1005 a_119_74# C1 a_32_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_386_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1007 a_32_74# B1 a_386_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_340_390# B2 a_27_390# VPB pshort w=1e+06u l=180000u
+  ad=6.8e+11p pd=5.36e+06u as=0p ps=0u
M1009 a_27_390# C2 a_32_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_390# B1 a_340_390# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_340_390# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.686e+11p ps=5.71e+06u
M1012 VPWR A2 a_340_390# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_32_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a222o_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
M1000 a_557_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.795e+11p pd=3.77e+06u as=9.428e+11p ps=7.49e+06u
M1001 a_119_392# C1 a_27_82# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=5.6e+11p ps=5.12e+06u
M1002 a_27_82# C2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_642_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=9.035e+11p pd=6.05e+06u as=1.10505e+12p ps=8.89e+06u
M1004 a_114_82# C1 a_27_82# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=4.832e+11p ps=4.07e+06u
M1005 X a_27_82# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 X a_27_82# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1007 a_27_82# A1 a_557_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_27_82# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_642_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_27_82# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_775_74# B1 a_27_82# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1012 VGND B2 a_775_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_392# B1 a_642_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_642_368# B2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND C2 a_114_82# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
M1000 VGND C2 a_119_74# VNB nlowvt w=640000u l=150000u
+  ad=9.312e+11p pd=5.47e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_119_392# C1 Y VPB pshort w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=6.1e+11p ps=5.22e+06u
M1002 a_461_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1003 a_119_74# C1 Y VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.92e+11p ps=4.41e+06u
M1004 Y B1 a_461_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_697_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1006 a_697_74# A1 Y VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_369_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.8e+11p pd=7.76e+06u as=4.2e+11p ps=2.84e+06u
M1008 VPWR A1 a_369_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_392# B2 a_369_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_369_392# B1 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a222oi_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
M1000 VGND A2 a_981_74# VNB nlowvt w=640000u l=150000u
+  ad=1.01862e+12p pd=8.5e+06u as=4.032e+11p ps=3.82e+06u
M1001 a_981_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_119_392# C2 Y VPB pshort w=1e+06u l=180000u
+  ad=1.17e+12p pd=1.034e+07u as=9.1e+11p ps=7.82e+06u
M1003 Y C1 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_137_74# C1 Y VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=7.232e+11p ps=7.38e+06u
M1005 a_981_74# A1 Y VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_981_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_119_392# B1 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.37e+12p ps=1.274e+07u
M1008 VGND C2 a_137_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B2 a_593_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1010 a_137_74# C2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C1 a_137_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_515_392# B2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_392# B2 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_515_392# B1 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_593_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_119_392# C1 Y VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=5.7e+11p pd=5.14e+06u as=0p ps=0u
M1018 Y C2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_515_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_593_74# B1 Y VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A2 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_515_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y B1 a_593_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_225_392# B1 a_230_79# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.344e+11p ps=1.7e+06u
M1001 VGND A2 a_52_123# VNB nlowvt w=640000u l=150000u
+  ad=4.426e+11p pd=4.38e+06u as=3.52e+11p ps=3.66e+06u
M1002 X a_225_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=8.412e+11p ps=5.86e+06u
M1003 a_230_79# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_135_392# B1 a_225_392# VPB pshort w=1e+06u l=180000u
+  ad=6.3e+11p pd=5.26e+06u as=3e+11p ps=2.6e+06u
M1005 a_135_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_225_392# B2 a_135_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_52_123# A1 a_225_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_225_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1009 VPWR A1 a_135_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_391_368# B2 a_81_48# VPB pshort w=1e+06u l=180000u
+  ad=6.1e+11p pd=5.22e+06u as=3.2e+11p ps=2.64e+06u
M1001 VPWR A2 a_391_368# VPB pshort w=1e+06u l=180000u
+  ad=9.412e+11p pd=8.24e+06u as=0p ps=0u
M1002 VGND a_81_48# X VNB nlowvt w=740000u l=150000u
+  ad=6.808e+11p pd=6.28e+06u as=2.072e+11p ps=2.04e+06u
M1003 a_81_48# B1 a_391_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_304_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=0p ps=0u
M1005 X a_81_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 a_491_74# B1 a_81_48# VNB nlowvt w=740000u l=150000u
+  ad=1.85e+11p pd=1.98e+06u as=2.59e+11p ps=2.18e+06u
M1007 VPWR a_81_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_81_48# A1 a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_81_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_391_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B2 a_491_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_645_120# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.89825e+11p pd=3.8e+06u as=1.217e+12p ps=1.055e+07u
M1001 a_95_306# B1 a_645_120# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1002 a_1064_123# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1003 a_95_306# A1 a_1064_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_555_392# VPB pshort w=1e+06u l=180000u
+  ad=1.6398e+12p pd=1.381e+07u as=1.36e+12p ps=1.272e+07u
M1005 X a_95_306# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1006 a_555_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_95_306# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_95_306# B2 a_555_392# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1009 X a_95_306# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1010 VPWR a_95_306# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_95_306# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_555_392# B1 a_95_306# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1064_123# A1 a_95_306# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_95_306# B1 a_555_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_95_306# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A2 a_555_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_95_306# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_645_120# B1 a_95_306# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_555_392# B2 a_95_306# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_95_306# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_555_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B2 a_645_120# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A2 a_1064_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_159_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1001 a_159_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.922e+11p ps=4.02e+06u
M1002 VPWR A1 a_71_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=9.184e+11p ps=8.36e+06u
M1003 a_339_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1004 Y B2 a_71_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 a_71_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_71_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_339_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_66_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.4896e+12p pd=1.386e+07u as=9.52e+11p ps=6.18e+06u
M1001 a_148_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=4.662e+11p ps=4.22e+06u
M1002 Y A1 a_148_74# VNB nlowvt w=740000u l=150000u
+  ad=7.918e+11p pd=6.58e+06u as=0p ps=0u
M1003 Y B1 a_66_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.384e+11p pd=5.62e+06u as=0p ps=0u
M1004 VGND A2 a_148_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_558_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.958e+11p pd=4.3e+06u as=0p ps=0u
M1006 Y B1 a_558_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B2 a_558_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_66_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_66_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_66_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_66_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B2 a_66_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_148_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_558_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_66_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_45_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.6992e+12p pd=2.498e+07u as=1.4672e+12p ps=1.158e+07u
M1001 a_48_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.0138e+12p pd=1.014e+07u as=8.288e+11p ps=8.16e+06u
M1002 a_48_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B2 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=0p ps=0u
M1004 a_45_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B2 a_48_74# VNB nlowvt w=740000u l=150000u
+  ad=8.288e+11p pd=8.16e+06u as=0p ps=0u
M1006 Y B2 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_45_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_840_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.0138e+12p pd=1.014e+07u as=0p ps=0u
M1010 a_48_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_45_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_840_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_840_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_48_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_840_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B1 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A1 a_840_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_45_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_45_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A1 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A2 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_45_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_45_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B1 a_48_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B1 a_48_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A2 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A1 a_840_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND B2 a_48_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_840_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_840_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A1 a_45_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR a_93_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=6.662e+11p pd=5.51e+06u as=2.912e+11p ps=2.76e+06u
M1001 a_261_392# A1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1002 a_93_264# a_257_126# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=8.3095e+11p ps=6.71e+06u
M1003 a_605_126# B2 a_93_264# VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1004 a_257_126# A1_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=0p ps=0u
M1005 VGND A2_N a_257_126# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_93_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1007 a_257_126# A2_N a_261_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1008 VGND B1 a_605_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_533_392# a_257_126# a_93_264# VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=2.6e+11p ps=2.52e+06u
M1010 a_533_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B2 a_533_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 X a_221_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=9.212e+11p ps=8.2e+06u
M1001 X a_221_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.184e+12p ps=9.5e+06u
M1002 VPWR a_221_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_221_74# B2 a_149_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1004 a_293_333# A2_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=0p ps=0u
M1005 VPWR B1 a_61_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.3e+11p ps=5.06e+06u
M1006 VGND a_293_333# a_221_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_149_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_221_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_61_392# B2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1_N a_549_378# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1011 VGND A1_N a_293_333# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_221_74# a_293_333# a_61_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1013 a_549_378# A2_N a_293_333# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VGND a_162_48# X VNB nlowvt w=740000u l=150000u
+  ad=1.6403e+12p pd=1.199e+07u as=4.144e+11p ps=4.08e+06u
M1001 a_1009_74# B2 a_162_48# VNB nlowvt w=640000u l=150000u
+  ad=5.184e+11p pd=5.46e+06u as=3.753e+11p ps=3.85e+06u
M1002 a_586_368# A1_N VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.352e+11p pd=2.66e+06u as=1.5368e+12p ps=1.358e+07u
M1003 a_162_48# a_586_94# a_820_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.06e+12p ps=1.012e+07u
M1004 a_820_392# a_586_94# a_162_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1009_74# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_586_94# A2_N a_586_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1007 X a_162_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 a_1009_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B2 a_820_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_162_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_162_48# B2 a_1009_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_162_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1013 a_820_392# B2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_586_94# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1015 VPWR B1 a_820_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_162_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_162_48# a_586_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_162_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_820_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_162_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_162_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2_N a_586_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_126_112# A1_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=8.322e+11p ps=6.72e+06u
M1001 Y a_126_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1002 a_126_112# A2_N a_120_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1003 VGND B1 a_488_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1004 a_402_368# a_126_112# Y VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=2.912e+11p ps=2.76e+06u
M1005 a_402_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.96e+11p ps=5.36e+06u
M1006 VPWR B2 a_402_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_488_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_120_392# A1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2_N a_126_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_615_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=5.994e+11p ps=6.06e+06u
M1001 a_212_392# A1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=8.648e+11p ps=8.08e+06u
M1002 Y a_212_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.17e+11p ps=8.02e+06u
M1003 Y a_212_102# a_424_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1872e+12p ps=1.108e+07u
M1004 a_424_368# a_212_102# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_615_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_615_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2_N a_212_102# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.93e+06u
M1008 VPWR B2 a_424_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_424_368# B2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_424_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_212_102# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_212_102# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_424_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B1 a_615_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_212_102# A2_N a_212_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_914_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0138e+12p pd=1.014e+07u as=1.2654e+12p ps=1.23e+07u
M1001 Y B2 a_914_74# VNB nlowvt w=740000u l=150000u
+  ad=8.288e+11p pd=8.16e+06u as=0p ps=0u
M1002 a_539_368# B2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.0944e+12p pd=1.942e+07u as=1.4796e+12p ps=1.366e+07u
M1003 VGND a_117_392# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_117_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B2 a_539_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1_N a_117_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1007 a_539_368# B2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B1 a_539_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B2 a_914_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_539_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1 a_914_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_914_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_914_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_117_392# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_117_392# a_539_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1016 VPWR B1 a_539_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_117_392# A2_N a_29_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u
M1018 a_29_392# A2_N a_117_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_539_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A1_N a_29_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_539_368# a_117_392# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_29_392# A1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_117_392# a_539_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_539_368# a_117_392# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND B1 a_914_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR B2 a_539_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_117_392# A2_N VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_117_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_914_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_261_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=8.9e+11p ps=5.96e+06u
M1001 VGND B1 a_89_270# VNB nlowvt w=640000u l=150000u
+  ad=5.289e+11p pd=4.33e+06u as=3.488e+11p ps=3.65e+06u
M1002 VPWR A2 a_261_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_89_270# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_264_120# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=2.10625e+11p pd=1.96e+06u as=0p ps=0u
M1005 a_89_270# C1 a_549_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1006 VGND a_89_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1007 a_89_270# A1 a_359_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1008 a_261_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_549_392# B1 a_261_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_89_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1011 a_359_123# A2 a_264_120# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR a_21_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.1724e+12p pd=8.7e+06u as=3.024e+11p ps=2.78e+06u
M1001 a_423_74# A2 a_351_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1002 VGND a_21_270# X VNB nlowvt w=740000u l=150000u
+  ad=7.955e+11p pd=6.59e+06u as=2.072e+11p ps=2.04e+06u
M1003 a_663_392# B1 a_333_392# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=6e+11p ps=5.2e+06u
M1004 VGND B1 a_21_270# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.847e+11p ps=4.27e+06u
M1005 a_351_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_21_270# C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_21_270# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2 a_333_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_333_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_333_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_21_270# A1 a_423_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_21_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_21_270# C1 a_663_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_157_392# C1 a_69_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u
M1001 a_69_392# C1 a_157_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND B1 a_157_392# VNB nlowvt w=640000u l=150000u
+  ad=1.23862e+12p pd=1.191e+07u as=5.376e+11p ps=5.52e+06u
M1003 VGND a_157_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1004 VPWR A3 a_337_392# VPB pshort w=1e+06u l=180000u
+  ad=1.7898e+12p pd=1.611e+07u as=1.08e+12p ps=1.016e+07u
M1005 a_337_392# B1 a_69_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_337_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_157_392# A1 a_1081_39# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=6.927e+11p ps=6.48e+06u
M1008 a_337_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1081_39# A1 a_157_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_337_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_337_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_69_392# B1 a_337_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_157_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_888_105# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1015 a_1081_39# A2 a_888_105# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A3 a_888_105# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND C1 a_157_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_157_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_157_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1020 a_888_105# A2 a_1081_39# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_157_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_157_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_157_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_157_392# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_157_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_337_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_157_392# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_159_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=7.952e+11p ps=5.9e+06u
M1001 a_231_74# A2 a_159_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1002 Y C1 a_465_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=3.36e+11p ps=2.84e+06u
M1003 a_465_368# B1 a_159_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=4.847e+11p ps=4.27e+06u
M1005 a_159_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_159_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2 a_159_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=7.178e+11p ps=4.9e+06u
M1001 a_130_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=1.2208e+12p ps=1.114e+07u
M1002 a_130_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A2 a_130_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_130_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_130_368# B1 a_692_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=8.848e+11p ps=8.3e+06u
M1006 a_692_368# B1 a_130_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C1 a_692_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1008 a_45_74# A2 a_300_74# VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=4.144e+11p ps=4.08e+06u
M1009 a_45_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A3 a_45_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A1 a_300_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_692_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_300_74# A2 a_45_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_300_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_130_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A3 a_130_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_117_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.4192e+12p pd=2.224e+07u as=2.0944e+12p ps=1.942e+07u
M1001 a_117_368# B1 a_1213_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.512e+12p ps=1.39e+07u
M1002 a_465_74# A2 a_34_74# VNB nlowvt w=740000u l=150000u
+  ad=8.288e+11p pd=8.16e+06u as=1.0286e+12p ps=1.018e+07u
M1003 a_34_74# A2 a_465_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A1 a_465_74# VNB nlowvt w=740000u l=150000u
+  ad=1.0286e+12p pd=1.018e+07u as=0p ps=0u
M1005 VPWR A2 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1213_368# B1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_465_74# A2 a_34_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_117_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C1 a_1213_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1010 VGND A3 a_34_74# VNB nlowvt w=740000u l=150000u
+  ad=1.4578e+12p pd=9.86e+06u as=0p ps=0u
M1011 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A2 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1213_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y C1 a_1213_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_465_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_117_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_34_74# A2 a_465_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A1 a_465_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1213_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A3 a_34_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_465_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_34_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_34_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_117_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A3 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_117_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_117_368# B1 a_1213_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR A3 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1213_368# B1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VGND B1 a_81_270# VNB nlowvt w=640000u l=150000u
+  ad=5.827e+11p pd=4.47e+06u as=2.816e+11p ps=2.16e+06u
M1001 a_253_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=9.8e+11p ps=6.14e+06u
M1002 a_81_270# B1 a_253_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1003 a_253_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A2 a_253_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_337_120# A2 a_265_120# VNB nlowvt w=640000u l=150000u
+  ad=2.5125e+11p pd=2.09e+06u as=1.344e+11p ps=1.7e+06u
M1006 VGND a_81_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1007 VPWR a_81_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1008 a_265_120# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_81_270# A1 a_337_120# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VGND B1 a_97_296# VNB nlowvt w=740000u l=150000u
+  ad=9.435e+11p pd=6.99e+06u as=3.108e+11p ps=2.32e+06u
M1001 a_371_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1002 X a_97_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.3546e+12p ps=9.02e+06u
M1003 VPWR a_97_296# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_365_368# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1005 VPWR A2 a_365_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_449_74# A2 a_371_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1007 VGND a_97_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1008 X a_97_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_365_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_97_296# B1 a_365_368# VPB pshort w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1011 a_97_296# A1 a_449_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_529_392# VPB pshort w=1e+06u l=180000u
+  ad=2.1676e+12p pd=1.682e+07u as=1.57e+12p ps=1.314e+07u
M1001 X a_83_274# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1002 a_83_274# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=5.888e+11p pd=5.68e+06u as=1.0507e+12p ps=1.001e+07u
M1003 VGND A3 a_1000_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.44e+11p ps=5.54e+06u
M1004 VPWR A2 a_529_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_83_274# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_775_74# A2 a_1000_74# VNB nlowvt w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=0p ps=0u
M1007 VGND B1 a_83_274# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_274# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_83_274# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_83_274# B1 a_529_392# VPB pshort w=1e+06u l=180000u
+  ad=3.4e+11p pd=2.68e+06u as=0p ps=0u
M1011 a_529_392# B1 a_83_274# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_83_274# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1013 VGND a_83_274# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_83_274# A1 a_775_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_775_74# A1 a_83_274# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1000_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1000_74# A2 a_775_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_83_274# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_83_274# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_529_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A3 a_529_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_529_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_529_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VPWR A2 a_139_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=6.14e+06u as=6.608e+11p ps=5.66e+06u
M1001 a_139_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B1 a_139_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1003 Y A1 a_223_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=3.108e+11p ps=2.32e+06u
M1004 a_223_74# A2 a_145_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1005 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.291e+11p pd=4.39e+06u as=0p ps=0u
M1006 a_145_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_139_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_200_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=7.548e+11p ps=5e+06u
M1001 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.217e+11p ps=4.37e+06u
M1002 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.6464e+12p pd=1.414e+07u as=9.744e+11p ps=8.46e+06u
M1003 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A1 a_200_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A3 a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1007 a_114_74# A2 a_200_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1010 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_114_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_200_74# A2 a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 Y A1 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=9.2695e+11p pd=8.48e+06u as=1.1544e+12p ps=9.04e+06u
M1001 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.272e+11p pd=5.6e+06u as=3.4272e+12p ps=2.628e+07u
M1002 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.0944e+12p ps=1.718e+07u
M1003 a_475_74# A2 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.03482e+12p ps=1.022e+07u
M1004 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_475_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_30_74# A2 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_30_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.2839e+12p ps=7.91e+06u
M1016 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A3 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_30_74# A2 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_475_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A1 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_475_74# A2 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A3 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_30_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_247_368# B2 a_84_48# VPB pshort w=1e+06u l=180000u
+  ad=8.2e+11p pd=7.64e+06u as=3.7e+11p ps=2.74e+06u
M1001 a_247_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.0496e+12p ps=6.26e+06u
M1002 a_84_48# B1 a_247_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_247_368# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A2 a_247_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_601_94# B1 a_84_48# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=4.032e+11p ps=2.54e+06u
M1006 a_259_94# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=6.004e+11p ps=4.48e+06u
M1007 a_337_94# A2 a_259_94# VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1008 VPWR a_84_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1009 VGND B2 a_601_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_84_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 a_84_48# A1 a_337_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_349_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.2e+11p pd=7.64e+06u as=1.417e+12p ps=9.14e+06u
M1001 a_45_264# B1 a_349_368# VPB pshort w=1e+06u l=180000u
+  ad=3.7e+11p pd=2.74e+06u as=0p ps=0u
M1002 a_661_74# B1 a_45_264# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=3.108e+11p ps=2.32e+06u
M1003 VGND a_45_264# X VNB nlowvt w=740000u l=150000u
+  ad=8.769e+11p pd=6.81e+06u as=2.146e+11p ps=2.06e+06u
M1004 X a_45_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VPWR a_45_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_433_74# A2 a_355_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=1.776e+11p ps=1.96e+06u
M1007 a_355_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B2 a_661_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_45_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_349_368# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_45_264# A1 a_433_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A2 a_349_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_349_368# B2 a_45_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_587_110# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=1.47252e+12p ps=1.141e+07u
M1001 a_83_283# B1 a_587_110# VNB nlowvt w=640000u l=150000u
+  ad=4.34975e+11p pd=4.13e+06u as=0p ps=0u
M1002 a_992_122# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=5.568e+11p pd=5.58e+06u as=0p ps=0u
M1003 X a_83_283# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=2.0706e+12p ps=1.665e+07u
M1004 X a_83_283# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_83_283# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_83_283# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_283# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=4.11e+06u as=0p ps=0u
M1008 X a_83_283# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_992_122# A2 a_1079_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.096e+11p ps=3.84e+06u
M1010 VPWR A2 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.955e+12p ps=1.591e+07u
M1011 a_509_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A3 a_992_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_509_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_83_283# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_509_392# B2 a_83_283# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.4e+11p ps=5.28e+06u
M1016 a_509_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A3 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_509_392# B1 a_83_283# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_83_283# B1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_83_283# B2 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_587_110# B1 a_83_283# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B2 a_587_110# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_83_283# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1079_122# A2 a_992_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_83_283# A1 a_1079_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1079_122# A1 a_83_283# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_119_74# VNB nlowvt w=740000u l=150000u
+  ad=6.068e+11p pd=3.12e+06u as=1.776e+11p ps=1.96e+06u
M1001 VGND A3 a_469_74# VNB nlowvt w=740000u l=150000u
+  ad=4.403e+11p pd=4.15e+06u as=3.108e+11p ps=2.32e+06u
M1002 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.0976e+12p pd=8.68e+06u as=3.584e+11p ps=2.88e+06u
M1003 Y B2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=9.968e+11p ps=6.26e+06u
M1005 a_119_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_391_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1009 a_469_74# A2 a_391_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=7.112e+11p pd=5.75e+06u as=2.1504e+12p ps=1.728e+07u
M1001 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.5288e+12p pd=9.45e+06u as=0p ps=0u
M1003 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_771_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.995e+11p pd=4.31e+06u as=6.66e+11p ps=6.24e+06u
M1006 a_27_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=6.808e+11p ps=6.28e+06u
M1008 Y A1 a_507_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=6.475e+11p ps=6.19e+06u
M1009 VGND A3 a_771_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_507_74# A2 a_771_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_771_74# A2 a_507_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_507_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.372e+12p pd=1.141e+07u as=3.8024e+12p ps=3.143e+07u
M1001 a_868_74# A2 a_1313_74# VNB nlowvt w=740000u l=150000u
+  ad=1.0471e+12p pd=1.023e+07u as=8.288e+11p ps=8.16e+06u
M1002 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.3128e+12p pd=1.757e+07u as=0p ps=0u
M1003 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A3 a_1313_74# VNB nlowvt w=740000u l=150000u
+  ad=1.1433e+12p pd=1.049e+07u as=0p ps=0u
M1005 a_868_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.806e+11p ps=8.3e+06u
M1006 a_1313_74# A2 a_868_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0952e+12p pd=1.036e+07u as=0p ps=0u
M1009 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1313_74# A2 a_868_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_868_74# A2 a_1313_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A3 a_1313_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_868_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y A1 a_868_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y A1 a_868_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1313_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1313_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_543_74# A2 a_449_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=2.368e+11p ps=2.12e+06u
M1001 VPWR a_83_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.1036e+12p pd=8.38e+06u as=3.136e+11p ps=2.8e+06u
M1002 a_357_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1003 a_449_74# A1 a_83_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 VPWR A3 a_357_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_83_244# X VNB nlowvt w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=7.104e+11p ps=3.4e+06u
M1006 a_657_74# A3 a_543_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1007 a_357_392# A4 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_83_244# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A4 a_657_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_357_392# B1 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1011 VPWR A1 a_357_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR a_441_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.6592e+12p pd=1.164e+07u as=3.024e+11p ps=2.78e+06u
M1001 a_441_74# B1 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=8.2e+11p ps=7.64e+06u
M1002 VPWR A4 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B1 a_441_74# VNB nlowvt w=740000u l=150000u
+  ad=1.1063e+12p pd=7.43e+06u as=2.886e+11p ps=2.26e+06u
M1004 a_199_74# A3 a_121_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=1.776e+11p ps=1.96e+06u
M1005 a_121_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_313_74# A2 a_199_74# VNB nlowvt w=740000u l=150000u
+  ad=3.626e+11p pd=2.46e+06u as=0p ps=0u
M1007 a_441_74# A1 a_313_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_441_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.034e+11p pd=2.3e+06u as=0p ps=0u
M1010 VPWR A2 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_441_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_441_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_113_98# B1 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=1.885e+12p ps=1.577e+07u
M1001 VGND a_113_98# X VNB nlowvt w=740000u l=150000u
+  ad=1.5409e+12p pd=1.26e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_1205_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1003 a_1205_74# A3 a_1010_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1004 X a_113_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_751_74# A2 a_1010_74# VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1006 a_113_98# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 a_27_392# A4 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.451e+12p ps=1.943e+07u
M1008 a_27_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A3 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A4 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_113_98# A1 a_751_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_751_74# A1 a_113_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A4 a_1205_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_113_98# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 a_113_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1010_74# A3 a_1205_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_113_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1022 VPWR a_113_98# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_113_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_113_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_113_98# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1010_74# A2 a_751_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_392# B1 a_113_98# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 VPWR A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1648e+12p pd=6.56e+06u as=9.744e+11p ps=8.46e+06u
M1001 Y A1 a_469_74# VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=3.108e+11p ps=2.32e+06u
M1002 VPWR A4 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_119_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1004 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_277_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=4.921e+11p ps=2.81e+06u
M1006 a_355_74# A3 a_277_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1007 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_469_74# A2 a_355_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.016e+12p pd=1.704e+07u as=1.7584e+12p ps=1.21e+07u
M1001 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_709_74# A3 a_512_74# VNB nlowvt w=740000u l=150000u
+  ad=6.438e+11p pd=6.18e+06u as=4.144e+11p ps=4.08e+06u
M1005 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=2.88e+06u
M1008 VPWR A4 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_239_74# A2 a_512_74# VNB nlowvt w=740000u l=150000u
+  ad=6.808e+11p pd=6.28e+06u as=0p ps=0u
M1011 Y A1 a_239_74# VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=0p ps=0u
M1012 a_27_368# A4 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.069e+11p ps=4.33e+06u
M1014 a_709_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A4 a_709_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_512_74# A2 a_239_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_512_74# A3 a_709_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_239_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.4664e+12p pd=3.083e+07u as=2.828e+12p ps=2.297e+07u
M1001 VPWR A4 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.552e+11p pd=5.65e+06u as=0p ps=0u
M1003 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1235_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0434e+12p pd=1.022e+07u as=8.658e+11p ps=8.26e+06u
M1005 a_852_74# A2 a_325_74# VNB nlowvt w=740000u l=150000u
+  ad=8.806e+11p pd=8.3e+06u as=1.3468e+12p ps=1.104e+07u
M1006 a_325_74# A2 a_852_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1235_74# A3 a_852_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_368# A4 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=7.252e+11p ps=6.4e+06u
M1016 VGND A4 a_1235_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A4 a_1235_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_852_74# A3 a_1235_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A1 a_325_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_852_74# A3 a_1235_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_325_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_325_74# A2 a_852_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A1 a_325_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_852_74# A2 a_325_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1235_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A4 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1235_74# A3 a_852_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_325_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_27_368# A4 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2_1 A B VGND VNB VPB VPWR X
M1000 a_56_136# A VPWR VPB pshort w=840000u l=180000u
+  ad=2.688e+11p pd=2.32e+06u as=6.076e+11p ps=5.2e+06u
M1001 VPWR B a_56_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_56_136# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1003 VGND B a_143_136# VNB nlowvt w=640000u l=150000u
+  ad=3.107e+11p pd=2.34e+06u as=2.752e+11p ps=2.28e+06u
M1004 a_143_136# A a_56_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1005 X a_56_136# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2_2 A B VGND VNB VPB VPWR X
M1000 VPWR B a_31_74# VPB pshort w=1e+06u l=180000u
+  ad=9.324e+11p pd=8.22e+06u as=2.7e+11p ps=2.54e+06u
M1001 X a_31_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1002 a_31_74# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B a_118_74# VNB nlowvt w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=1.776e+11p ps=1.96e+06u
M1004 VPWR a_31_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_31_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 a_118_74# A a_31_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1007 VGND a_31_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2_4 A B VGND VNB VPB VPWR X
M1000 VGND a_83_269# X VNB nlowvt w=740000u l=150000u
+  ad=8.594e+11p pd=8.14e+06u as=5.254e+11p ps=4.38e+06u
M1001 X a_83_269# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_83_269# A a_504_119# VNB nlowvt w=640000u l=150000u
+  ad=2.08e+11p pd=1.93e+06u as=3.872e+11p ps=3.77e+06u
M1003 VGND a_83_269# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_504_119# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_504_119# A a_83_269# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_83_269# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.272e+11p pd=5.6e+06u as=1.46945e+12p ps=1.304e+07u
M1007 VPWR a_83_269# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B a_504_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_83_269# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_83_269# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A a_83_269# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.746e+11p ps=4.49e+06u
M1012 X a_83_269# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_83_269# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_83_269# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B a_83_269# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2b_1 A_N B VGND VNB VPB VPWR X
M1000 VGND B a_353_98# VNB nlowvt w=640000u l=150000u
+  ad=6.2665e+11p pd=4.56e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_353_98# a_27_74# a_266_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1002 X a_266_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=6.594e+11p ps=5.27e+06u
M1003 X a_266_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=8.4e+11p ps=3.68e+06u
M1005 a_266_98# a_27_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1006 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1007 VPWR B a_266_98# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2b_2 A_N B VGND VNB VPB VPWR X
M1000 a_505_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=8.742e+11p ps=5.41e+06u
M1001 a_198_48# a_27_74# a_505_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1002 VPWR a_198_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.45745e+12p pd=9.24e+06u as=3.024e+11p ps=2.78e+06u
M1003 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1004 VGND a_198_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 a_198_48# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1006 VPWR a_27_74# a_198_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1008 X a_198_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_198_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2b_4 A_N B VGND VNB VPB VPWR X
M1000 VPWR B a_221_424# VPB pshort w=840000u l=180000u
+  ad=1.574e+12p pd=1.352e+07u as=4.536e+11p ps=4.44e+06u
M1001 VGND a_221_424# X VNB nlowvt w=740000u l=150000u
+  ad=9.074e+11p pd=8.29e+06u as=4.218e+11p ps=4.1e+06u
M1002 X a_221_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1003 VPWR a_221_424# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_221_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_221_424# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_221_424# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_221_424# a_27_392# a_233_74# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=4.16e+11p ps=3.86e+06u
M1008 VPWR A_N a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1009 a_233_74# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1011 X a_221_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_221_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_233_74# a_27_392# a_221_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_221_424# a_27_392# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B a_233_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_392# a_221_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_221_424# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3_1 A B C VGND VNB VPB VPWR X
M1000 X a_27_398# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.00785e+12p ps=6.04e+06u
M1001 a_121_136# A a_27_398# VNB nlowvt w=640000u l=150000u
+  ad=2.624e+11p pd=2.1e+06u as=1.824e+11p ps=1.85e+06u
M1002 a_233_136# B a_121_136# VNB nlowvt w=640000u l=150000u
+  ad=2.22e+11p pd=2.09e+06u as=0p ps=0u
M1003 a_27_398# B VPWR VPB pshort w=840000u l=180000u
+  ad=4.62e+11p pd=4.46e+06u as=0p ps=0u
M1004 VGND C a_233_136# VNB nlowvt w=640000u l=150000u
+  ad=3.107e+11p pd=2.34e+06u as=0p ps=0u
M1005 VPWR C a_27_398# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_27_398# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_398# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3_2 A B C VGND VNB VPB VPWR X
M1000 X a_41_384# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=6.9565e+11p ps=5.12e+06u
M1001 X a_41_384# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.2592e+12p ps=8.72e+06u
M1002 VPWR a_41_384# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND C a_247_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1004 a_247_136# B a_133_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.12e+06u
M1005 a_133_136# A a_41_384# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1006 VPWR A a_41_384# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.62e+11p ps=4.46e+06u
M1007 a_41_384# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C a_41_384# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_41_384# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3_4 A B C VGND VNB VPB VPWR X
M1000 a_686_74# B a_489_74# VNB nlowvt w=640000u l=150000u
+  ad=5.76e+11p pd=5.64e+06u as=3.84e+11p ps=3.76e+06u
M1001 VPWR B a_83_260# VPB pshort w=840000u l=180000u
+  ad=2.184e+12p pd=1.636e+07u as=7.14e+11p ps=6.74e+06u
M1002 a_489_74# B a_686_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1004 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_83_260# C VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C a_83_260# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_489_74# C VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=9.013e+11p ps=8.26e+06u
M1010 a_83_260# A a_686_74# VNB nlowvt w=640000u l=150000u
+  ad=2.368e+11p pd=2.02e+06u as=0p ps=0u
M1011 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1012 a_83_260# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_83_260# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C a_489_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_83_260# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_686_74# A a_83_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3b_1 A_N B C VGND VNB VPB VPWR X
M1000 a_266_94# B VPWR VPB pshort w=840000u l=180000u
+  ad=4.662e+11p pd=4.47e+06u as=9.786e+11p ps=7.71e+06u
M1001 X a_266_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_114_74# A_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.73e+11p pd=2.33e+06u as=0p ps=0u
M1003 X a_266_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=5.5385e+11p ps=4.28e+06u
M1004 a_353_94# a_114_74# a_266_94# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.824e+11p ps=1.85e+06u
M1005 a_431_94# B a_353_94# VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1006 a_114_74# A_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.9525e+11p pd=1.81e+06u as=0p ps=0u
M1007 VGND C a_431_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C a_266_94# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_114_74# a_266_94# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3b_2 A_N B C VGND VNB VPB VPWR X
M1000 VGND C a_454_74# VNB nlowvt w=740000u l=150000u
+  ad=6.8395e+11p pd=6.06e+06u as=3.108e+11p ps=2.32e+06u
M1001 a_284_368# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.5e+11p pd=5.1e+06u as=1.3408e+12p ps=1.08e+07u
M1002 VPWR a_27_88# a_284_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR C a_284_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_284_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VPWR A_N a_27_88# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 a_454_74# B a_376_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1007 X a_284_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1008 a_376_74# a_27_88# a_284_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 VGND A_N a_27_88# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1010 VGND a_284_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_284_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3b_4 A_N B C VGND VNB VPB VPWR X
M1000 VPWR A_N a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=2.3986e+12p pd=1.727e+07u as=2.8e+11p ps=2.56e+06u
M1001 VPWR a_301_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.048e+11p ps=5.56e+06u
M1002 a_239_98# a_27_74# a_301_368# VNB nlowvt w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=1.792e+11p ps=1.84e+06u
M1003 a_498_98# C VGND VNB nlowvt w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=1.063e+12p ps=1.005e+07u
M1004 VGND a_301_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1005 a_301_368# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.1e+11p pd=7.62e+06u as=0p ps=0u
M1006 VPWR C a_301_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_301_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_301_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_498_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_239_98# B a_498_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_498_98# B a_239_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_301_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_301_368# a_27_74# a_239_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_301_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_301_368# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_301_368# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_301_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A_N a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1019 VPWR B a_301_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_27_74# a_301_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_301_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__buf_1 A VGND VNB VPB VPWR X
M1000 X a_27_164# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=3.808e+11p ps=2.98e+06u
M1001 VPWR A a_27_164# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1002 VGND A a_27_164# VNB nlowvt w=550000u l=150000u
+  ad=3.0395e+11p pd=2.34e+06u as=2.4915e+11p ps=2.37e+06u
M1003 X a_27_164# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4_1 A B C D VGND VNB VPB VPWR X
M1000 VPWR B a_96_74# VPB pshort w=840000u l=180000u
+  ad=1.1326e+12p pd=8.13e+06u as=5.376e+11p ps=4.64e+06u
M1001 VPWR D a_96_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_96_74# C VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND D a_335_74# VNB nlowvt w=640000u l=150000u
+  ad=2.554e+11p pd=2.2e+06u as=2.688e+11p ps=2.12e+06u
M1004 a_96_74# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_96_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 X a_96_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1007 a_257_74# B a_179_74# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.536e+11p ps=1.76e+06u
M1008 a_335_74# C a_257_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_179_74# A a_96_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4_2 A B C D VGND VNB VPB VPWR X
M1000 a_221_74# B a_143_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=1.776e+11p ps=1.96e+06u
M1001 a_56_74# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=1.7568e+12p ps=1.184e+07u
M1002 VGND a_56_74# X VNB nlowvt w=740000u l=150000u
+  ad=5.846e+11p pd=4.54e+06u as=2.072e+11p ps=2.04e+06u
M1003 VPWR B a_56_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND D a_335_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.108e+11p ps=2.32e+06u
M1005 a_143_74# A a_56_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1006 a_56_74# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR D a_56_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_56_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_56_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1010 VPWR a_56_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_335_74# C a_221_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4_4 A B C D VGND VNB VPB VPWR X
M1000 X a_119_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.608e+11p pd=5.66e+06u as=2.657e+12p ps=1.983e+07u
M1001 a_119_392# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.145e+12p pd=1.029e+07u as=0p ps=0u
M1002 VPWR A a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_119_392# A a_119_119# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=3.584e+11p ps=3.68e+06u
M1004 a_119_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_119_119# B a_32_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.321e+11p ps=5.54e+06u
M1006 a_119_119# A a_119_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_119_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_119_392# X VNB nlowvt w=740000u l=150000u
+  ad=1.05515e+12p pd=8.94e+06u as=4.366e+11p ps=4.14e+06u
M1009 X a_119_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_119_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_119_392# D VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_392# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR D a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND D a_463_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1017 X a_119_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_32_119# B a_119_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_463_119# C a_32_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_463_119# D VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_32_119# C a_463_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_119_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_119_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4b_1 A_N B C D VGND VNB VPB VPWR X
M1000 VGND D a_526_139# VNB nlowvt w=640000u l=150000u
+  ad=4.5645e+11p pd=3.97e+06u as=3.418e+11p ps=2.55e+06u
M1001 a_448_139# B a_353_124# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=2.21125e+11p ps=2.08e+06u
M1002 a_229_424# a_27_74# VPWR VPB pshort w=840000u l=180000u
+  ad=5.628e+11p pd=4.7e+06u as=1.5316e+12p ps=9.08e+06u
M1003 a_353_124# a_27_74# a_229_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1004 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1005 X a_229_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 VPWR B a_229_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1008 VPWR D a_229_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_229_424# C VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_229_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1011 a_526_139# C a_448_139# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4b_2 A_N B C D VGND VNB VPB VPWR X
M1000 a_459_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=7.2205e+11p ps=4.95e+06u
M1001 a_537_74# C a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1002 a_186_48# D VPWR VPB pshort w=1e+06u l=180000u
+  ad=6.05e+11p pd=5.21e+06u as=1.75605e+12p ps=1.211e+07u
M1003 a_186_48# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_186_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 VPWR A_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 VPWR C a_186_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_186_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1008 a_645_74# B a_537_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1009 VPWR a_186_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1011 VPWR a_27_112# a_186_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_186_48# a_27_112# a_645_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 X a_186_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4b_4 A_N B C D VGND VNB VPB VPWR X
M1000 a_664_125# C a_751_125# VNB nlowvt w=640000u l=150000u
+  ad=5.37125e+11p pd=5.53e+06u as=3.872e+11p ps=3.77e+06u
M1001 VPWR a_199_294# X VPB pshort w=1.12e+06u l=180000u
+  ad=2.605e+12p pd=1.972e+07u as=7.28e+11p ps=5.78e+06u
M1002 a_664_125# B a_1136_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.992e+11p ps=4.12e+06u
M1003 a_199_294# D VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.64e+12p pd=1.128e+07u as=0p ps=0u
M1004 VPWR A_N a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1005 VGND a_199_294# X VNB nlowvt w=740000u l=150000u
+  ad=1.25925e+12p pd=9.57e+06u as=4.144e+11p ps=4.08e+06u
M1006 a_199_294# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND D a_751_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_27_368# a_199_294# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_199_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_199_294# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A_N a_27_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1012 a_199_294# a_27_368# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1136_125# a_27_368# a_199_294# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1014 X a_199_294# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_199_294# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_751_125# C a_664_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_199_294# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B a_199_294# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1136_125# B a_664_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR D a_199_294# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_751_125# D VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_199_294# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_199_294# a_27_368# a_1136_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR C a_199_294# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_199_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
M1000 VGND D a_647_74# VNB nlowvt w=640000u l=150000u
+  ad=5.299e+11p pd=4.38e+06u as=2.304e+11p ps=2e+06u
M1001 X a_179_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1002 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=1.2502e+12p pd=1.007e+07u as=2.352e+11p ps=2.24e+06u
M1003 a_455_74# a_27_74# a_179_48# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.824e+11p ps=1.85e+06u
M1004 a_533_74# a_503_48# a_455_74# VNB nlowvt w=640000u l=150000u
+  ad=2.688e+11p pd=2.12e+06u as=0p ps=0u
M1005 a_179_48# C VPWR VPB pshort w=840000u l=180000u
+  ad=4.956e+11p pd=4.54e+06u as=0p ps=0u
M1006 VPWR D a_179_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_503_48# a_179_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_179_48# a_27_74# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_503_48# B_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1010 a_503_48# B_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1011 a_647_74# C a_533_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_179_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=4.648e+11p pd=3.07e+06u as=0p ps=0u
M1013 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_225_82# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.1e+11p pd=5.62e+06u as=1.854e+12p ps=1.212e+07u
M1001 VPWR D a_225_82# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_390_82# a_354_252# a_312_82# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.776e+11p ps=1.96e+06u
M1003 X a_225_82# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.0454e+12p ps=7.35e+06u
M1004 a_312_82# a_27_74# a_225_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1005 a_354_252# B_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1006 a_354_252# B_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1007 VGND a_225_82# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_225_82# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 VPWR a_225_82# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_498_82# C a_390_82# VNB nlowvt w=740000u l=150000u
+  ad=2.664e+11p pd=2.2e+06u as=0p ps=0u
M1011 VGND D a_498_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_354_252# a_225_82# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_225_82# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1015 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_685_140# a_27_74# a_412_140# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=5.888e+11p ps=5.68e+06u
M1001 a_685_140# C a_882_137# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.888e+11p ps=5.68e+06u
M1002 a_412_140# a_27_74# a_685_140# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR B_N a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=3.5296e+12p pd=2.358e+07u as=2.8e+11p ps=2.56e+06u
M1004 a_475_388# D VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.3525e+12p pd=1.087e+07u as=0p ps=0u
M1005 X a_475_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1006 VPWR a_475_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_475_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_475_388# X VNB nlowvt w=740000u l=150000u
+  ad=1.1064e+12p pd=1.017e+07u as=4.44e+11p ps=4.16e+06u
M1009 a_475_388# a_200_74# a_412_140# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1010 VGND D a_882_137# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_475_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_475_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_475_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR D a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_475_388# a_200_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_475_388# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_200_74# a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR C a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_27_74# a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_475_388# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_475_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_200_74# A_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1023 VGND B_N a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1024 a_200_74# A_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.915e+11p pd=1.99e+06u as=0p ps=0u
M1025 a_882_137# C a_685_140# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_882_137# D VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_412_140# a_200_74# a_475_388# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__buf_16 A VGND VNB VPB VPWR X
M1000 a_83_260# A VGND VNB nlowvt w=740000u l=150000u
+  ad=6.734e+11p pd=6.26e+06u as=2.8305e+12p ps=2.541e+07u
M1001 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.6576e+12p pd=1.632e+07u as=0p ps=0u
M1002 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A a_83_260# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=3.7632e+12p pd=3.36e+07u as=2.4192e+12p ps=2.224e+07u
M1005 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_83_260# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A a_83_260# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_83_260# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_83_260# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.072e+11p pd=8.34e+06u as=0p ps=0u
M1023 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A a_83_260# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_83_260# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A a_83_260# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_83_260# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR A a_83_260# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_83_260# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__buf_2 A VGND VNB VPB VPWR X
M1000 X a_21_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1278e+12p ps=6.51e+06u
M1001 VPWR a_21_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_21_260# X VNB nlowvt w=740000u l=150000u
+  ad=5.216e+11p pd=4.39e+06u as=2.072e+11p ps=2.04e+06u
M1003 a_21_260# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1004 a_21_260# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.05e+11p pd=2.61e+06u as=0p ps=0u
M1005 X a_21_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__buf_4 A VGND VNB VPB VPWR X
M1000 VGND a_86_260# X VNB nlowvt w=740000u l=150000u
+  ad=1.1063e+12p pd=7.43e+06u as=4.144e+11p ps=4.08e+06u
M1001 a_86_260# A VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=1.2278e+12p ps=1.077e+07u
M1002 VPWR A a_86_260# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_86_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_86_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_86_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.048e+11p ps=5.56e+06u
M1006 X a_86_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_86_260# A VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 X a_86_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_86_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_86_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__buf_8 A VGND VNB VPB VPWR X
M1000 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=8.325e+11p pd=8.17e+06u as=1.591e+12p ps=1.318e+07u
M1001 VPWR A a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=1.9768e+12p pd=1.697e+07u as=6.16e+11p ps=5.58e+06u
M1002 a_27_74# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.2824e+12p ps=1.125e+07u
M1005 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=0p ps=0u
M1007 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__bufbuf_16 A VGND VNB VPB VPWR X
M1000 a_588_74# a_203_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=3.3855e+12p ps=2.987e+07u
M1001 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.6576e+12p ps=1.632e+07u
M1002 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.4752e+12p pd=2.234e+07u as=4.3344e+12p ps=3.91e+07u
M1003 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_588_74# a_203_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.072e+11p pd=8.34e+06u as=0p ps=0u
M1005 VGND a_203_74# a_588_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_203_74# a_588_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1012 a_203_74# a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=0p ps=0u
M1013 a_588_74# a_203_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_588_74# a_203_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_27_368# a_203_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_203_74# a_588_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_203_74# a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_203_74# a_588_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_203_74# a_588_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_27_368# a_203_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.181e+11p ps=4.09e+06u
M1034 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_588_74# a_203_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_203_74# a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 X a_588_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_588_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_588_74# a_203_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_588_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 X a_588_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND a_203_74# a_588_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VGND A a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1051 a_203_74# a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__bufbuf_8 A VGND VNB VPB VPWR X
M1000 a_224_368# a_27_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=2.2302e+12p ps=1.971e+07u
M1001 VGND a_334_368# X VNB nlowvt w=740000u l=150000u
+  ad=1.7549e+12p pd=1.515e+07u as=8.732e+11p ps=8.28e+06u
M1002 VPWR a_334_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.2656e+12p ps=1.122e+07u
M1003 X a_334_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_334_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_334_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_334_368# a_224_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=0p ps=0u
M1007 X a_334_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_334_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_334_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_334_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1012 X a_334_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_334_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_224_368# a_27_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1015 VGND a_224_368# a_334_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1017 X a_334_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_224_368# a_334_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.16e+11p ps=5.58e+06u
M1019 VGND a_224_368# a_334_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_334_368# a_224_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_334_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_334_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_334_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_224_368# a_334_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_334_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__bufinv_16 A VGND VNB VPB VPWR Y
M1000 a_27_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=3.2079e+12p ps=2.791e+07u
M1001 VPWR A a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=4.0656e+12p pd=3.638e+07u as=6.16e+11p ps=5.58e+06u
M1002 a_27_74# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.6576e+12p ps=1.632e+07u
M1004 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.464e+12p pd=2.232e+07u as=0p ps=0u
M1005 VPWR A a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_384_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=8.38e+06u as=0p ps=0u
M1010 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_384_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1012 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_27_74# a_384_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_74# a_384_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_27_74# a_384_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_384_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_27_74# a_384_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_27_74# a_384_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_384_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_27_74# a_384_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Y a_384_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VGND a_384_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR a_384_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Y a_384_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_384_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_384_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__bufinv_8 A VGND VNB VPB VPWR Y
M1000 a_183_48# a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=1.9824e+12p ps=1.698e+07u
M1001 VPWR a_183_48# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.3552e+12p ps=1.138e+07u
M1002 Y a_183_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_183_48# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_27_368# a_183_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_183_48# a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_183_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=8.954e+11p pd=8.34e+06u as=1.5392e+12p ps=1.304e+07u
M1007 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 Y a_183_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_183_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_183_48# a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.292e+11p pd=4.12e+06u as=0p ps=0u
M1011 VPWR a_183_48# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_183_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_183_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_183_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_183_48# a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_183_48# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_183_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_183_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_27_368# a_183_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_183_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y a_183_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_183_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkbuf_1 A VGND VNB VPB VPWR X
M1000 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=4.144e+11p ps=2.98e+06u
M1001 VPWR A a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1002 X a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.19e+11p pd=1.41e+06u as=3.276e+11p ps=2.4e+06u
M1003 VGND A a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkbuf_16 A VGND VNB VPB VPWR X
M1000 a_114_74# A VGND VNB nlowvt w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=1.4826e+12p ps=1.63e+07u
M1001 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=9.408e+11p ps=1.12e+07u
M1002 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_114_74# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=3.3824e+12p ps=3.068e+07u
M1004 VPWR A a_114_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.4192e+12p pd=2.224e+07u as=0p ps=0u
M1006 a_114_74# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_114_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A a_114_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_114_74# A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND A a_114_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_114_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 X a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 X a_114_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_114_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkbuf_2 A VGND VNB VPB VPWR X
M1000 X a_43_192# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=6.048e+11p ps=5.56e+06u
M1001 VPWR a_43_192# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_43_192# A VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=2.667e+11p ps=2.95e+06u
M1003 a_43_192# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1004 X a_43_192# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1005 VGND a_43_192# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkbuf_4 A VGND VNB VPB VPWR X
M1000 VGND a_83_270# X VNB nlowvt w=420000u l=150000u
+  ad=3.969e+11p pd=4.41e+06u as=2.52e+11p ps=2.88e+06u
M1001 X a_83_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.744e+11p ps=8.46e+06u
M1002 VPWR a_83_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_83_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_83_270# A VGND VNB nlowvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1005 a_83_270# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1006 VPWR a_83_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_270# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_270# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_270# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkbuf_8 A VGND VNB VPB VPWR X
M1000 VGND a_128_74# X VNB nlowvt w=420000u l=150000u
+  ad=8.757e+11p pd=9.21e+06u as=4.809e+11p ps=5.65e+06u
M1001 VGND a_128_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_128_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2264e+12p pd=1.115e+07u as=2.0552e+12p ps=1.711e+07u
M1003 VPWR a_128_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A a_128_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1005 X a_128_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_128_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_128_74# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_128_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_128_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_128_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_128_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A a_128_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1013 X a_128_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_128_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_128_74# A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_128_74# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_128_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_128_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_128_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkdlyinv3sd1_1 A VGND VNB VPB VPWR Y
M1000 Y a_288_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=1.0312e+12p ps=6.42e+06u
M1001 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1002 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1003 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=4.2e+11p pd=3.68e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 Y a_288_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkdlyinv3sd2_1 A VGND VNB VPB VPWR Y
M1000 Y a_288_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=9.312e+11p ps=6.22e+06u
M1001 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=4.074e+11p ps=3.62e+06u
M1002 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1003 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=250000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1005 Y a_288_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkdlyinv3sd3_1 A VGND VNB VPB VPWR Y
M1000 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=500000u
+  ad=2.6e+11p pd=2.52e+06u as=6.812e+11p ps=5.72e+06u
M1001 Y a_288_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1002 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=4.074e+11p ps=3.62e+06u
M1003 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1004 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 Y a_288_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkdlyinv5sd1_1 A VGND VNB VPB VPWR Y
M1000 a_549_74# a_288_74# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.65e+11p pd=2.53e+06u as=1.8512e+12p ps=1.006e+07u
M1001 a_549_74# a_288_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=7.623e+11p ps=6.15e+06u
M1002 Y a_682_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 VPWR a_549_74# a_682_74# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=6.1e+11p ps=3.22e+06u
M1004 VGND a_549_74# a_682_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.583e+11p ps=2.07e+06u
M1005 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1006 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1007 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 Y a_682_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1009 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkdlyinv5sd2_1 A VGND VNB VPB VPWR Y
M1000 a_549_74# a_288_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=7.371e+11p ps=6.03e+06u
M1001 VGND a_549_74# a_682_74# VNB nlowvt w=420000u l=180000u
+  ad=0p pd=0u as=2.457e+11p ps=2.01e+06u
M1002 Y a_682_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 a_549_74# a_288_74# VPWR VPB pshort w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=1.6512e+12p ps=9.66e+06u
M1004 VPWR a_549_74# a_682_74# VPB pshort w=1e+06u l=250000u
+  ad=0p pd=0u as=5.1e+11p ps=3.02e+06u
M1005 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1007 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 Y a_682_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1009 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=250000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkdlyinv5sd3_1 A VGND VNB VPB VPWR Y
M1000 VPWR a_549_74# a_682_74# VPB pshort w=1e+06u l=500000u
+  ad=1.1512e+12p pd=8.66e+06u as=2.6e+11p ps=2.52e+06u
M1001 a_549_74# a_288_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=7.371e+11p ps=6.03e+06u
M1002 VGND a_549_74# a_682_74# VNB nlowvt w=420000u l=180000u
+  ad=0p pd=0u as=2.457e+11p ps=2.01e+06u
M1003 Y a_682_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1004 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=500000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1005 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1007 a_549_74# a_288_74# VPWR VPB pshort w=1e+06u l=500000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1008 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 Y a_682_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkinv_1 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=2.2535e+11p pd=2.17e+06u as=1.491e+11p ps=1.55e+06u
M1001 Y A VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u
M1002 VPWR A Y VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkinv_16 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.696e+12p pd=3.348e+07u as=4.0656e+12p ps=3.638e+07u
M1001 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=9.408e+11p pd=1.12e+07u as=1.83765e+12p ps=1.762e+07u
M1002 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkinv_2 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=6.16e+11p ps=5.58e+06u
M1001 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=2.394e+11p pd=2.82e+06u as=3.276e+11p ps=2.4e+06u
M1003 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkinv_4 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=4.242e+11p pd=3.7e+06u as=6.216e+11p ps=5.48e+06u
M1001 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.072e+11p pd=8.34e+06u as=1.344e+12p ps=1.136e+07u
M1003 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkinv_8 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=1.2264e+12p pd=9.2e+06u as=7.77e+11p ps=7.9e+06u
M1001 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.8144e+12p pd=1.668e+07u as=2.4472e+12p ps=2.005e+07u
M1003 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR short w=510000u l=45000u
R1 VGND LO short w=510000u l=45000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__decap_4 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB pshort w=1e+06u l=1e+06u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nlowvt w=420000u l=1e+06u
+  ad=2.31e+11p pd=2.78e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__decap_8 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB pshort w=1e+06u l=1e+06u
+  ad=8.35e+11p pd=7.67e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nlowvt w=420000u l=1e+06u
+  ad=3.465e+11p pd=4.17e+06u as=0p ps=0u
M1002 VPWR VGND VPWR VPB pshort w=1e+06u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND VPWR VGND VNB nlowvt w=420000u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 VGND a_1534_446# a_1611_140# VNB nlowvt w=420000u l=150000u
+  ad=1.55002e+12p pd=1.351e+07u as=1.008e+11p ps=1.32e+06u
M1001 a_595_119# a_27_74# a_523_119# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1002 VGND a_1534_446# a_2412_410# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 VPWR a_978_357# a_936_424# VPB pshort w=840000u l=180000u
+  ad=2.39652e+12p pd=2.021e+07u as=1.764e+11p ps=2.1e+06u
M1004 Q_N a_1534_446# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1005 a_311_119# a_200_74# a_595_119# VNB nlowvt w=420000u l=150000u
+  ad=5.1975e+11p pd=3.99e+06u as=0p ps=0u
M1006 a_540_503# a_474_405# VPWR VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 a_1300_424# a_474_405# VPWR VPB pshort w=840000u l=180000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1008 VGND RESET_B a_978_357# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1009 Q a_2412_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1010 a_523_119# a_474_405# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR RESET_B a_978_357# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1012 a_311_119# a_27_74# a_595_119# VPB pshort w=420000u l=180000u
+  ad=3.3585e+11p pd=3.41e+06u as=1.386e+11p ps=1.5e+06u
M1013 a_474_405# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=4.452e+11p pd=4.42e+06u as=0p ps=0u
M1014 VGND D a_311_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_595_119# a_200_74# a_540_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1818_76# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=5.032e+11p pd=4.56e+06u as=0p ps=0u
M1017 VPWR D a_311_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1486_508# a_27_74# a_1349_114# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.688e+11p ps=2.4e+06u
M1019 a_1920_392# a_978_357# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1020 a_474_405# a_595_119# a_867_119# VNB nlowvt w=550000u l=150000u
+  ad=1.925e+11p pd=1.8e+06u as=3.4925e+11p ps=3.47e+06u
M1021 a_936_424# a_595_119# a_474_405# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1611_140# a_200_74# a_1349_114# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=6.2825e+11p ps=3.42e+06u
M1023 VPWR a_1534_446# a_1486_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1254_119# a_474_405# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.83125e+11p pd=1.8e+06u as=0p ps=0u
M1025 VPWR SET_B a_1534_446# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.45e+11p ps=5.09e+06u
M1026 a_1534_446# a_1349_114# a_1920_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND SET_B a_867_119# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1349_114# a_27_74# a_1254_119# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q_N a_1534_446# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1030 VPWR CLK_N a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1031 a_200_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1032 a_867_119# a_978_357# a_474_405# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1818_76# a_1349_114# a_1534_446# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1034 a_1534_446# a_978_357# a_1818_76# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND CLK_N a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1036 a_200_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1037 Q a_2412_410# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1038 a_1349_114# a_200_74# a_1300_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_1534_446# a_2412_410# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1555_410# a_1335_112# a_1934_392# VPB pshort w=1e+06u l=180000u
+  ad=5.45e+11p pd=5.09e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR a_1555_410# a_2516_368# VPB pshort w=1e+06u l=180000u
+  ad=3.0275e+12p pd=2.579e+07u as=2.65e+11p ps=2.53e+06u
M1002 a_1507_508# a_27_74# a_1335_112# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.688e+11p ps=2.4e+06u
M1003 a_1240_125# a_473_405# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.90125e+11p pd=1.88e+06u as=2.06398e+12p ps=1.857e+07u
M1004 a_1640_138# a_200_74# a_1335_112# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=6.1e+11p ps=3.85e+06u
M1005 VGND SET_B a_867_125# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=3.4925e+11p ps=3.47e+06u
M1006 a_933_424# a_601_119# a_473_405# VPB pshort w=840000u l=180000u
+  ad=2.016e+11p pd=2.16e+06u as=4.452e+11p ps=4.42e+06u
M1007 a_867_125# a_975_322# a_473_405# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.54e+11p ps=1.66e+06u
M1008 Q a_2516_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1009 a_1832_74# a_1335_112# a_1555_410# VNB nlowvt w=740000u l=150000u
+  ad=4.979e+11p pd=4.43e+06u as=2.368e+11p ps=2.12e+06u
M1010 a_1832_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_311_119# a_27_74# a_601_119# VPB pshort w=420000u l=180000u
+  ad=3.3075e+11p pd=3.39e+06u as=1.386e+11p ps=1.5e+06u
M1012 VPWR RESET_B a_975_322# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1013 VPWR a_1555_410# a_1507_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_473_405# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q_N a_1555_410# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1016 Q a_2516_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1017 VGND D a_311_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=5.0085e+11p ps=3.93e+06u
M1018 a_539_503# a_473_405# VPWR VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1019 VPWR a_1555_410# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_2516_368# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1934_392# a_975_322# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1335_112# a_200_74# a_1315_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.016e+11p ps=2.16e+06u
M1023 VGND a_1555_410# a_1640_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1555_410# a_975_322# a_1832_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR D a_311_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND RESET_B a_975_322# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1027 VPWR SET_B a_1555_410# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_311_119# a_200_74# a_601_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1029 VPWR a_975_322# a_933_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_601_119# a_200_74# a_539_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_1555_410# a_2516_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1032 VGND a_2516_368# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR CLK_N a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1034 a_200_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1035 VGND a_1555_410# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1036 a_529_119# a_473_405# VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1037 VGND CLK_N a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1038 a_200_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1039 a_1335_112# a_27_74# a_1240_125# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_473_405# a_601_119# a_867_125# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1315_424# a_473_405# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_601_119# a_27_74# a_529_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Q_N a_1555_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR RESET_B a_1062_93# VPB pshort w=640000u l=180000u
+  ad=2.7277e+12p pd=2.199e+07u as=1.664e+11p ps=1.8e+06u
M1001 a_1421_508# a_214_74# a_1314_424# VPB pshort w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=2.667e+11p ps=2.39e+06u
M1002 Q_N a_1474_446# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.83492e+12p ps=1.558e+07u
M1003 a_1206_379# a_671_93# VPWR VPB pshort w=840000u l=180000u
+  ad=3.339e+11p pd=2.85e+06u as=0p ps=0u
M1004 a_520_87# a_27_74# a_422_125# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.7605e+11p ps=1.9e+06u
M1005 a_1314_424# a_27_74# a_1206_379# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1318_119# a_671_93# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1007 VGND RESET_B a_1062_93# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1008 Q_N a_1474_446# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1009 VPWR a_671_93# a_716_379# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 a_1817_392# a_1314_424# a_1474_446# VPB pshort w=1e+06u l=180000u
+  ad=2.35e+11p pd=2.47e+06u as=3.35e+11p ps=2.67e+06u
M1011 VPWR a_1062_93# a_1020_379# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.016e+11p ps=2.16e+06u
M1012 a_1314_424# a_214_74# a_1318_119# VNB nlowvt w=550000u l=150000u
+  ad=2.317e+11p pd=2.33e+06u as=0p ps=0u
M1013 a_422_125# D VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1014 a_1498_74# a_27_74# a_1314_424# VNB nlowvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1015 VPWR a_1474_446# a_1421_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_520_87# a_214_74# a_422_125# VPB pshort w=420000u l=180000u
+  ad=2.163e+11p pd=2.36e+06u as=0p ps=0u
M1017 a_214_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1018 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1019 VGND a_1474_446# a_2320_410# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1020 a_671_93# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=3.024e+11p pd=2.4e+06u as=0p ps=0u
M1021 VGND a_1474_446# a_1498_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_671_93# a_520_87# a_872_119# VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=6.465e+11p ps=4.96e+06u
M1023 a_1474_446# SET_B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1062_93# a_1817_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_606_87# a_214_74# a_520_87# VNB nlowvt w=420000u l=150000u
+  ad=1.645e+11p pd=1.81e+06u as=0p ps=0u
M1026 VPWR a_1474_446# a_2320_410# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1027 a_1474_446# a_1314_424# a_1708_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=4.884e+11p ps=4.28e+06u
M1028 a_214_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1029 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1030 a_872_119# a_1062_93# a_671_93# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1708_74# a_1062_93# a_1474_446# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_422_125# D VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_872_119# SET_B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1708_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1020_379# a_520_87# a_671_93# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_671_93# a_606_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q a_2320_410# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1038 Q a_2320_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1039 a_716_379# a_27_74# a_520_87# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1434_74# a_307_387# a_1224_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=4.33e+11p ps=3.08e+06u
M1001 a_910_119# a_841_401# a_832_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1002 a_841_401# a_709_463# VGND VNB nlowvt w=640000u l=150000u
+  ad=3.222e+11p pd=2.44e+06u as=1.3521e+12p ps=1.212e+07u
M1003 a_1224_74# a_501_387# a_841_401# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Q a_2026_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_709_463# a_501_387# a_38_78# VPB pshort w=420000u l=180000u
+  ad=2.247e+11p pd=2.75e+06u as=2.31e+11p ps=2.78e+06u
M1006 VPWR CLK a_307_387# VPB pshort w=1.12e+06u l=180000u
+  ad=1.90045e+12p pd=1.771e+07u as=3.361e+11p ps=2.92e+06u
M1007 VPWR a_1482_48# a_1468_471# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 Q_N a_1224_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.72e+11p pd=3.44e+06u as=0p ps=0u
M1009 a_799_463# a_307_387# a_709_463# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 a_125_78# D a_38_78# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.394e+11p ps=2.82e+06u
M1011 VGND CLK a_307_387# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.45475e+11p ps=2.15e+06u
M1012 a_501_387# a_307_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.262e+11p pd=2.14e+06u as=0p ps=0u
M1013 VGND a_1224_74# a_2026_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1014 a_501_387# a_307_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 Q_N a_1224_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1016 a_841_401# a_709_463# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1017 a_832_119# a_501_387# a_709_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1018 a_709_463# a_307_387# a_38_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND RESET_B a_910_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1224_74# a_307_387# a_841_401# VPB pshort w=1e+06u l=180000u
+  ad=3.664e+11p pd=3.14e+06u as=0p ps=0u
M1021 a_1482_48# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1022 VGND a_1482_48# a_1434_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_38_78# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR RESET_B a_38_78# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1224_74# a_1482_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1624_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1027 a_1482_48# a_1224_74# a_1624_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1028 VPWR a_841_401# a_799_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND RESET_B a_125_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1224_74# a_2026_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1031 a_709_463# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_2026_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1033 a_1468_471# a_501_387# a_1224_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 Q a_2366_352# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=3.6099e+12p ps=2.652e+07u
M1001 Q a_2366_352# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.19475e+12p ps=1.777e+07u
M1002 a_1800_291# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1003 VPWR a_2366_352# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR RESET_B a_70_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.864e+11p ps=3.52e+06u
M1005 a_1758_389# a_818_418# a_1586_149# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=3.55e+11p ps=3e+06u
M1006 a_298_294# a_728_331# a_70_74# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.632e+11p ps=3.03e+06u
M1007 a_728_331# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 VGND a_1800_291# a_1499_149# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1009 a_728_331# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1010 VGND a_1586_149# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1011 VPWR RESET_B a_298_294# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.247e+11p ps=2.75e+06u
M1012 a_156_74# D a_70_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 a_686_485# a_334_119# VPWR VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1014 VPWR a_1800_291# a_1758_389# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_614_81# a_334_119# a_536_81# VNB nlowvt w=420000u l=150000u
+  ad=3.465e+11p pd=3.33e+06u as=1.008e+11p ps=1.32e+06u
M1016 VGND a_2366_352# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1586_149# a_728_331# a_1499_149# VNB nlowvt w=420000u l=150000u
+  ad=2.165e+11p pd=2.13e+06u as=0p ps=0u
M1018 a_1800_291# a_1586_149# a_1974_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1019 VPWR a_1586_149# a_1800_291# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_2366_352# a_1586_149# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.75e+11p pd=2.75e+06u as=0p ps=0u
M1021 a_1974_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_2366_352# a_1586_149# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1023 a_334_119# a_298_294# VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.45e+11p pd=5.09e+06u as=0p ps=0u
M1024 a_298_294# a_728_331# a_686_485# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_334_119# a_818_418# a_1586_149# VNB nlowvt w=740000u l=150000u
+  ad=5.2345e+11p pd=4.67e+06u as=0p ps=0u
M1026 a_70_74# a_818_418# a_298_294# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1586_149# a_728_331# a_334_119# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_536_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_728_331# a_818_418# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.998e+11p ps=2.02e+06u
M1030 Q_N a_1586_149# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1031 a_334_119# a_298_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_614_81# a_818_418# a_298_294# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q_N a_1586_149# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_728_331# a_818_418# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1035 VPWR a_1586_149# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_70_74# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND RESET_B a_156_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
M1000 a_856_294# a_714_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.5e+11p pd=3.5e+06u as=1.65038e+12p ps=1.553e+07u
M1001 a_1266_119# a_510_74# a_856_294# VPB pshort w=1e+06u l=180000u
+  ad=4.264e+11p pd=3.34e+06u as=0p ps=0u
M1002 VGND a_1598_93# a_1550_119# VNB nlowvt w=420000u l=150000u
+  ad=1.2824e+12p pd=1.089e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_510_74# a_300_347# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1004 a_1598_93# a_1266_119# a_1736_119# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1005 VPWR a_856_294# a_820_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_714_119# a_510_74# a_33_74# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=2.31e+11p ps=2.78e+06u
M1007 a_1266_119# a_300_347# a_856_294# VNB nlowvt w=740000u l=150000u
+  ad=6.134e+11p pd=4.02e+06u as=2.146e+11p ps=2.06e+06u
M1008 VPWR a_1598_93# a_1550_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 VGND RESET_B a_922_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 a_1736_119# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_510_74# a_300_347# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.257e+11p pd=2.09e+06u as=0p ps=0u
M1012 a_714_119# a_300_347# a_33_74# VPB pshort w=420000u l=180000u
+  ad=2.226e+11p pd=2.74e+06u as=2.31e+11p ps=2.78e+06u
M1013 VGND CLK_N a_300_347# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.442e+11p ps=2.14e+06u
M1014 a_820_457# a_510_74# a_714_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1598_93# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1016 a_922_119# a_856_294# a_850_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 VPWR CLK_N a_300_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9575e+11p ps=2.65e+06u
M1018 a_714_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_850_119# a_300_347# a_714_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_856_294# a_714_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1266_119# a_1934_94# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1022 a_1550_119# a_510_74# a_1266_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_1266_119# a_1598_93# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND RESET_B a_120_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VPWR a_1266_119# a_1934_94# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1026 Q a_1934_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 Q a_1934_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=0p ps=0u
M1028 a_120_74# D a_33_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1550_508# a_300_347# a_1266_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_33_74# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR RESET_B a_33_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_1656_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.33593e+12p ps=1.182e+07u
M1001 a_493_387# a_299_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.262e+11p pd=2.14e+06u as=0p ps=0u
M1002 a_821_138# a_493_387# a_701_463# VNB nlowvt w=420000u l=150000u
+  ad=9.03e+10p pd=1.27e+06u as=1.407e+11p ps=1.51e+06u
M1003 VGND a_1867_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 a_1266_74# a_299_387# a_833_400# VPB pshort w=1e+06u l=180000u
+  ad=4.39e+11p pd=3.4e+06u as=3.5125e+11p ps=2.95e+06u
M1005 VPWR a_1867_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=1.82245e+12p pd=1.716e+07u as=3.64e+11p ps=2.89e+06u
M1006 VGND RESET_B a_894_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_701_463# a_299_387# a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.541e+11p ps=2.89e+06u
M1008 VPWR a_833_400# a_791_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 VGND RESET_B a_117_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 a_1471_493# a_493_387# a_1266_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1011 a_1867_409# a_1266_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1012 a_894_138# a_833_400# a_821_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_1518_203# a_1476_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1014 a_701_463# a_493_387# a_30_78# VPB pshort w=420000u l=180000u
+  ad=2.31e+11p pd=2.78e+06u as=2.31e+11p ps=2.78e+06u
M1015 VPWR a_1518_203# a_1471_493# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1476_81# a_299_387# a_1266_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.58e+11p ps=3.28e+06u
M1017 a_1518_203# a_1266_74# a_1656_81# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1018 a_30_78# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR RESET_B a_30_78# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1518_203# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1021 VPWR CLK a_299_387# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.1375e+11p ps=2.92e+06u
M1022 a_791_463# a_299_387# a_701_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK a_299_387# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.45475e+11p ps=2.15e+06u
M1024 VPWR a_1266_74# a_1518_203# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_493_387# a_299_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1026 a_117_78# D a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1266_74# a_493_387# a_833_400# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.921e+11p ps=2.81e+06u
M1028 a_1867_409# a_1266_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1029 a_833_400# a_701_463# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_701_463# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_833_400# a_701_463# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_837_359# a_699_463# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.38125e+11p pd=2.8e+06u as=2.1627e+12p ps=1.993e+07u
M1001 VGND RESET_B a_895_138# VNB nlowvt w=420000u l=150000u
+  ad=1.91777e+12p pd=1.512e+07u as=1.008e+11p ps=1.32e+06u
M1002 VPWR a_1271_74# a_1525_212# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.226e+11p ps=1.9e+06u
M1003 a_1271_74# a_493_387# a_837_359# VNB nlowvt w=740000u l=150000u
+  ad=4.58e+11p pd=3.28e+06u as=2.405e+11p ps=2.13e+06u
M1004 a_699_463# a_493_387# a_30_78# VPB pshort w=420000u l=180000u
+  ad=2.31e+11p pd=2.78e+06u as=2.289e+11p ps=2.77e+06u
M1005 VGND a_1525_212# a_1481_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_789_463# a_306_119# a_699_463# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 a_1271_74# a_306_119# a_837_359# VPB pshort w=1e+06u l=180000u
+  ad=4.32625e+11p pd=3.6e+06u as=0p ps=0u
M1008 a_895_138# a_837_359# a_817_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 a_1481_493# a_493_387# a_1271_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1010 a_1924_409# a_1271_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1011 VPWR a_837_359# a_789_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND RESET_B a_117_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_493_387# a_306_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.98825e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_30_78# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR RESET_B a_30_78# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND CLK a_306_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_699_463# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1525_212# a_1481_493# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1525_212# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1924_409# a_1271_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_1663_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1022 a_1525_212# a_1271_74# a_1663_81# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1023 a_837_359# a_699_463# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_817_138# a_493_387# a_699_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1025 VPWR CLK a_306_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1026 a_699_463# a_306_119# a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.82e+06u
M1027 a_493_387# a_306_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1028 a_117_78# D a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q a_1924_409# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1030 VPWR a_1924_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Q a_1924_409# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1032 a_1481_81# a_306_119# a_1271_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_1924_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_702_463# a_303_395# a_37_78# VNB nlowvt w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=2.31e+11p ps=2.78e+06u
M1001 VGND CLK a_303_395# VNB nlowvt w=740000u l=150000u
+  ad=2.086e+12p pd=1.709e+07u as=2.45475e+11p ps=2.15e+06u
M1002 a_497_395# a_303_395# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.262e+11p pd=2.14e+06u as=0p ps=0u
M1003 VGND a_2013_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.847e+11p ps=4.27e+06u
M1004 a_1353_392# a_497_395# a_834_355# VNB nlowvt w=740000u l=150000u
+  ad=4.58e+11p pd=3.28e+06u as=9.435e+11p ps=4.03e+06u
M1005 VGND RESET_B a_124_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VPWR a_834_355# a_792_463# VPB pshort w=420000u l=180000u
+  ad=2.9869e+12p pd=2.378e+07u as=8.82e+10p ps=1.26e+06u
M1007 a_1630_493# a_497_395# a_1353_392# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=6.511e+11p ps=4.41e+06u
M1008 VPWR a_1353_392# a_2013_409# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1009 Q a_2013_409# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.552e+11p pd=5.65e+06u as=0p ps=0u
M1010 VPWR CLK a_303_395# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.32375e+11p ps=2.92e+06u
M1011 a_834_355# a_702_463# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_1678_395# a_1630_493# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_497_395# a_303_395# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1014 a_702_463# a_497_395# a_37_78# VPB pshort w=420000u l=180000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1015 a_834_355# a_702_463# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1016 a_702_463# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_124_78# D a_37_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_2013_409# a_1353_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 a_792_463# a_303_395# a_702_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1353_392# a_303_395# a_834_355# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_2013_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1678_395# a_1647_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1023 VGND a_2013_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_890_138# a_834_355# a_812_138# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1025 a_2013_409# a_1353_392# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1678_395# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1027 VPWR a_1353_392# a_1678_395# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Q a_2013_409# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2013_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1827_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1031 a_1678_395# a_1353_392# a_1827_81# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1032 Q a_2013_409# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND RESET_B a_890_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_37_78# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR RESET_B a_37_78# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_812_138# a_497_395# a_702_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1647_81# a_303_395# a_1353_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q a_2013_409# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1262_74# a_596_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=2.176e+11p pd=1.96e+06u as=1.56945e+12p ps=1.386e+07u
M1001 a_1257_341# a_596_81# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.565e+11p pd=3.01e+06u as=1.91615e+12p ps=1.7e+07u
M1002 a_1358_377# a_225_74# a_1257_341# VPB pshort w=1e+06u l=180000u
+  ad=5.371e+11p pd=4.81e+06u as=0p ps=0u
M1003 VGND D a_27_80# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.82e+06u
M1004 a_596_81# a_225_74# a_27_80# VNB nlowvt w=420000u l=150000u
+  ad=2.562e+11p pd=2.06e+06u as=0p ps=0u
M1005 a_1520_508# a_398_74# a_1358_377# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1006 VGND a_779_380# a_748_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_731_463# a_225_74# a_596_81# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.344e+11p ps=1.48e+06u
M1008 Q_N a_1358_377# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 a_596_81# a_398_74# a_27_80# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1010 VPWR a_1510_48# a_1520_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1510_48# a_1358_377# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1012 VPWR CLK a_225_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1013 a_398_74# a_225_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_1358_377# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1061_74# a_596_81# a_779_380# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.113e+11p ps=1.37e+06u
M1016 VPWR SET_B a_779_380# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1017 VPWR a_1358_377# a_1510_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.533e+11p ps=1.57e+06u
M1018 a_1358_377# a_398_74# a_1262_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1019 a_398_74# a_225_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1020 VPWR a_779_380# a_731_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q a_2113_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_748_81# a_398_74# a_596_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR D a_27_80# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND SET_B a_1540_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VGND a_1358_377# a_2113_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1026 VGND SET_B a_1061_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q a_2113_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1028 a_1540_74# a_1510_48# a_1462_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1029 a_779_380# a_596_81# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q_N a_1358_377# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1031 a_1462_74# a_225_74# a_1358_377# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND CLK a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1033 VPWR a_1358_377# a_2113_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR SET_B a_757_401# VPB pshort w=420000u l=180000u
+  ad=2.75e+12p pd=2.354e+07u as=1.407e+11p ps=1.51e+06u
M1001 a_595_97# a_398_74# a_27_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=2.352e+11p ps=2.8e+06u
M1002 VGND SET_B a_1531_118# VNB nlowvt w=420000u l=150000u
+  ad=2.28115e+12p pd=1.92e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_1501_92# a_1339_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
M1004 VGND a_2221_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 a_709_463# a_225_74# a_595_97# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1006 a_1261_341# a_595_97# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.69625e+11p pd=3.16e+06u as=0p ps=0u
M1007 VGND a_1339_74# a_2221_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1008 Q_N a_1339_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 VPWR a_757_401# a_709_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1524_508# a_398_74# a_1339_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=5.425e+11p ps=4.65e+06u
M1011 Q a_2221_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1012 a_1261_74# a_595_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1013 Q_N a_1339_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1014 VPWR a_2221_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_1339_74# a_2221_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1016 Q a_2221_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_595_97# a_225_74# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=2.394e+11p ps=2.82e+06u
M1018 VPWR CLK a_225_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1019 a_398_74# a_225_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1020 a_757_401# a_595_97# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_398_74# a_225_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1022 a_1339_74# a_398_74# a_1261_74# VNB nlowvt w=640000u l=150000u
+  ad=2.314e+11p pd=2.12e+06u as=0p ps=0u
M1023 a_1531_118# a_1501_92# a_1453_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1024 VGND a_1339_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_757_401# a_731_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1026 VPWR a_1339_74# a_1501_92# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.481e+11p ps=2.24e+06u
M1027 a_1339_74# a_225_74# a_1261_341# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND SET_B a_1001_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1029 VPWR D a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1339_74# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_1501_92# a_1524_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1001_74# a_595_97# a_757_401# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 VGND D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1339_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND CLK a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1036 a_731_97# a_398_74# a_595_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1453_118# a_225_74# a_1339_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
M1000 a_760_395# a_604_74# VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=1.7201e+12p ps=1.561e+07u
M1001 a_1200_341# a_604_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.69625e+11p pd=3.16e+06u as=0p ps=0u
M1002 VPWR a_1470_48# a_1460_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1003 a_1215_74# a_604_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=2.4e+11p pd=2.03e+06u as=1.40335e+12p ps=1.213e+07u
M1004 VPWR CLK a_224_350# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1005 a_1470_48# a_1301_392# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1006 a_1301_392# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=5.212e+11p pd=4.59e+06u as=0p ps=0u
M1007 a_1301_392# a_398_74# a_1215_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1008 VPWR D a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.31e+11p ps=2.78e+06u
M1009 VGND SET_B a_1027_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 a_398_74# a_224_350# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1011 a_1027_118# a_604_74# a_760_395# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1012 VPWR SET_B a_760_395# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_604_74# a_224_350# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=2.9565e+11p ps=3.17e+06u
M1014 Q a_1902_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1015 a_712_463# a_224_350# a_604_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.344e+11p ps=1.48e+06u
M1016 a_1470_48# a_1301_392# VPWR VPB pshort w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1017 a_604_74# a_398_74# a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1422_74# a_224_350# a_1301_392# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1019 a_1500_74# a_1470_48# a_1422_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1020 a_398_74# a_224_350# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1021 a_1301_392# a_224_350# a_1200_341# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_760_395# a_740_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1023 VGND SET_B a_1500_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_740_74# a_398_74# a_604_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_1902_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1026 VGND a_1301_392# a_1902_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1027 a_1460_508# a_398_74# a_1301_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1301_392# a_1902_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1030 VPWR a_760_395# a_712_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND CLK a_224_350# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
M1000 a_1278_74# a_612_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.6502e+12p ps=1.426e+07u
M1001 a_1356_74# a_398_74# a_1278_74# VNB nlowvt w=640000u l=150000u
+  ad=2.713e+11p pd=2.31e+06u as=0p ps=0u
M1002 a_1057_118# a_612_74# a_767_384# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1003 a_1356_74# a_225_74# a_1269_341# VPB pshort w=1e+06u l=180000u
+  ad=5.278e+11p pd=4.58e+06u as=3.69625e+11p ps=3.16e+06u
M1004 VGND SET_B a_1596_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1005 VGND a_2022_94# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1006 VPWR a_1356_74# a_2022_94# VPB pshort w=1e+06u l=180000u
+  ad=2.34017e+12p pd=1.968e+07u as=2.8e+11p ps=2.56e+06u
M1007 a_1356_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1489_118# a_225_74# a_1356_74# VNB nlowvt w=420000u l=150000u
+  ad=1.617e+11p pd=1.61e+06u as=0p ps=0u
M1009 a_767_384# a_612_74# VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1010 a_1524_508# a_398_74# a_1356_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1011 a_1269_341# a_612_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_781_74# a_398_74# a_612_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.919e+11p ps=2.23e+06u
M1013 VGND a_1356_74# a_2022_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1014 VPWR CLK a_225_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1015 a_398_74# a_225_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 VPWR SET_B a_767_384# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_398_74# a_225_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1018 a_612_74# a_225_74# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.0635e+11p ps=3.21e+06u
M1019 a_1566_92# a_1356_74# VPWR VPB pshort w=420000u l=180000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1020 VPWR D a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1021 a_719_456# a_225_74# a_612_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.344e+11p ps=1.48e+06u
M1022 VGND SET_B a_1057_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_612_74# a_398_74# a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_767_384# a_781_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_2022_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_2022_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 a_1566_92# a_1356_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1028 VPWR a_1566_92# a_1524_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2022_94# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1596_118# a_1566_92# a_1489_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_767_384# a_719_456# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND CLK a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
M1000 VGND a_1324_392# a_1940_74# VNB nlowvt w=740000u l=150000u
+  ad=2.1906e+12p pd=1.727e+07u as=2.627e+11p ps=2.19e+06u
M1001 a_612_74# a_398_74# a_27_74# VPB pshort w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=2.352e+11p ps=2.8e+06u
M1002 a_719_463# a_225_74# a_612_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1003 VGND a_767_402# a_732_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 VGND SET_B a_1514_88# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 a_1484_62# a_1324_392# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1006 a_1324_392# a_398_74# a_1225_74# VNB nlowvt w=640000u l=150000u
+  ad=2.1145e+11p pd=2e+06u as=2.528e+11p ps=2.07e+06u
M1007 a_1514_88# a_1484_62# a_1436_88# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 Q a_1940_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.477e+11p pd=4.17e+06u as=0p ps=0u
M1009 VGND a_1940_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_767_402# a_719_463# VPB pshort w=420000u l=180000u
+  ad=2.5187e+12p pd=2.304e+07u as=0p ps=0u
M1011 VPWR SET_B a_767_402# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1012 a_1484_62# a_1324_392# VPWR VPB pshort w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1013 a_732_74# a_398_74# a_612_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.89e+11p ps=1.74e+06u
M1014 VPWR a_1484_62# a_1483_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1015 a_1436_88# a_225_74# a_1324_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND SET_B a_1035_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1017 VGND a_1940_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_398_74# a_225_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 a_1324_392# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=5.212e+11p pd=4.59e+06u as=0p ps=0u
M1020 a_1940_74# a_1324_392# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1021 VPWR a_1324_392# a_1940_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q a_1940_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1023 a_612_74# a_225_74# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.0635e+11p ps=3.21e+06u
M1024 VPWR CLK a_225_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1025 a_1324_392# a_225_74# a_1223_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.64375e+11p ps=3.1e+06u
M1026 a_1035_118# a_612_74# a_767_402# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.491e+11p ps=1.55e+06u
M1027 a_398_74# a_225_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1028 a_1225_74# a_612_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1940_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q a_1940_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR D a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1223_347# a_612_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q a_1940_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND CLK a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1036 a_1483_508# a_398_74# a_1324_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_1940_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_767_402# a_612_74# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
M1000 Q_N a_1644_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=1.78195e+12p ps=1.538e+07u
M1001 VPWR a_1005_120# a_1191_120# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1002 a_546_447# a_27_74# a_423_503# VNB nlowvt w=420000u l=150000u
+  ad=1.51375e+11p pd=1.66e+06u as=1.176e+11p ps=1.4e+06u
M1003 a_653_508# a_27_74# a_546_447# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.02475e+11p ps=2.16e+06u
M1004 VPWR a_1191_120# a_1161_482# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 VGND a_701_463# a_713_102# VNB nlowvt w=420000u l=150000u
+  ad=1.71272e+12p pd=1.365e+07u as=8.82e+10p ps=1.26e+06u
M1006 Q a_1191_120# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VPWR a_1191_120# a_1644_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1008 a_701_463# a_546_447# VGND VNB nlowvt w=550000u l=150000u
+  ad=2.365e+11p pd=2.26e+06u as=0p ps=0u
M1009 a_423_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1005_120# a_208_368# a_701_463# VNB nlowvt w=550000u l=150000u
+  ad=2.593e+11p pd=2.18e+06u as=0p ps=0u
M1011 a_701_463# a_546_447# VPWR VPB pshort w=840000u l=180000u
+  ad=4.83e+11p pd=2.83e+06u as=0p ps=0u
M1012 a_713_102# a_208_368# a_546_447# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_1191_120# a_1143_146# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1014 a_208_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1015 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1016 a_1161_482# a_208_368# a_1005_120# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.628e+11p ps=2.39e+06u
M1017 a_208_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.252e+11p pd=2.59e+06u as=0p ps=0u
M1018 VGND a_1005_120# a_1191_120# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1019 VPWR a_701_463# a_653_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1143_146# a_27_74# a_1005_120# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_423_503# D VPWR VPB pshort w=420000u l=180000u
+  ad=2.8015e+11p pd=2.61e+06u as=0p ps=0u
M1022 VGND a_1191_120# a_1644_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1023 a_1005_120# a_27_74# a_701_463# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q a_1191_120# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1025 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 a_546_447# a_208_368# a_423_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_1644_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
M1000 a_1248_128# a_27_74# a_1003_424# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.9205e+11p ps=3.36e+06u
M1001 Q a_1290_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.10485e+12p ps=1.739e+07u
M1002 VGND a_753_284# a_717_102# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1003 Q_N a_1835_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 a_454_503# D VPWR VPB pshort w=420000u l=180000u
+  ad=1.9985e+11p pd=2.13e+06u as=2.66788e+12p ps=2.211e+07u
M1005 a_753_284# a_561_445# VGND VNB nlowvt w=550000u l=150000u
+  ad=3.87e+11p pd=2.98e+06u as=0p ps=0u
M1006 VGND a_1835_368# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_1835_368# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1008 a_1290_102# a_1003_424# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1009 VGND a_1290_102# a_1248_128# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1011 a_209_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1012 a_705_445# a_27_74# a_561_445# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.268e+11p ps=1.92e+06u
M1013 a_209_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.252e+11p pd=2.59e+06u as=0p ps=0u
M1014 a_753_284# a_561_445# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1015 a_1003_424# a_27_74# a_753_284# VPB pshort w=840000u l=180000u
+  ad=4.662e+11p pd=3.4e+06u as=0p ps=0u
M1016 VPWR a_1290_102# a_1835_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1017 VPWR a_1003_424# a_1290_102# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1003_424# a_209_368# a_753_284# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_1290_102# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_717_102# a_209_368# a_561_445# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.66075e+11p ps=1.73e+06u
M1021 VGND a_1290_102# a_1835_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1022 Q a_1290_102# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1023 VPWR a_1290_102# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_561_445# a_209_368# a_454_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1211_479# a_209_368# a_1003_424# VPB pshort w=420000u l=180000u
+  ad=1.659e+11p pd=1.63e+06u as=0p ps=0u
M1026 VPWR a_1290_102# a_1211_479# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_1835_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_1003_424# a_1290_102# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1029 VPWR a_753_284# a_705_445# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_454_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1031 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1032 a_561_445# a_27_74# a_454_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfxtp_1 CLK D VGND VNB VPB VPWR Q
M1000 VPWR a_1014_424# a_1210_314# VPB pshort w=840000u l=180000u
+  ad=1.41472e+12p pd=1.248e+07u as=2.352e+11p ps=2.24e+06u
M1001 a_1168_124# a_27_74# a_1014_424# VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.362e+11p ps=2.07e+06u
M1002 a_209_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.553e+11p pd=2.17e+06u as=1.2645e+12p ps=1.059e+07u
M1003 a_1014_424# a_27_74# a_713_458# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=4.41e+11p ps=2.73e+06u
M1004 a_713_458# a_564_463# VGND VNB nlowvt w=550000u l=150000u
+  ad=2.18125e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_1121_508# a_209_368# a_1014_424# VPB pshort w=420000u l=180000u
+  ad=1.869e+11p pd=1.73e+06u as=0p ps=0u
M1006 a_1014_424# a_209_368# a_713_458# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_457_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=3.1125e+11p pd=2.43e+06u as=0p ps=0u
M1008 VGND a_1014_424# a_1210_314# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1010 a_209_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1011 VPWR a_713_458# a_671_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 a_564_463# a_209_368# a_457_503# VPB pshort w=420000u l=180000u
+  ad=1.841e+11p pd=1.95e+06u as=1.841e+11p ps=1.95e+06u
M1013 Q a_1210_314# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 VGND a_713_458# a_731_101# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1015 a_671_503# a_27_74# a_564_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_731_101# a_209_368# a_564_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.575e+11p ps=1.73e+06u
M1017 a_564_463# a_27_74# a_457_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_713_458# a_564_463# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Q a_1210_314# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1020 a_457_503# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1210_314# a_1168_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 VPWR a_1210_314# a_1121_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfxtp_2 CLK D VGND VNB VPB VPWR Q
M1000 VGND a_695_459# a_708_101# VNB nlowvt w=420000u l=150000u
+  ad=1.65997e+12p pd=1.34e+07u as=1.008e+11p ps=1.32e+06u
M1001 VGND a_1217_314# a_1172_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1002 VPWR a_695_459# a_647_504# VPB pshort w=420000u l=180000u
+  ad=1.72835e+12p pd=1.511e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_695_459# a_541_429# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=0p ps=0u
M1004 a_695_459# a_541_429# VPWR VPB pshort w=840000u l=180000u
+  ad=4.998e+11p pd=2.87e+06u as=0p ps=0u
M1005 Q a_1217_314# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1217_314# a_1128_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.869e+11p ps=1.73e+06u
M1007 a_434_508# D VPWR VPB pshort w=420000u l=180000u
+  ad=2.18225e+11p pd=2.34e+06u as=0p ps=0u
M1008 Q a_1217_314# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 a_1022_424# a_209_368# a_695_459# VNB nlowvt w=550000u l=150000u
+  ad=2.4555e+11p pd=2.35e+06u as=0p ps=0u
M1010 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1011 a_209_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1012 a_541_429# a_209_368# a_434_508# VPB pshort w=420000u l=180000u
+  ad=2.12625e+11p pd=2.29e+06u as=0p ps=0u
M1013 a_434_508# D VGND VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1014 VPWR a_1217_314# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_708_101# a_209_368# a_541_429# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.5225e+11p ps=1.67e+06u
M1016 a_541_429# a_27_74# a_434_508# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1172_124# a_27_74# a_1022_424# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1022_424# a_27_74# a_695_459# VPB pshort w=840000u l=180000u
+  ad=2.625e+11p pd=2.38e+06u as=0p ps=0u
M1019 VPWR a_1022_424# a_1217_314# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1020 VGND a_1022_424# a_1217_314# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1021 VGND a_1217_314# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_647_504# a_27_74# a_541_429# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1128_508# a_209_368# a_1022_424# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1025 a_209_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.775e+11p pd=2.23e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfxtp_4 CLK D VGND VNB VPB VPWR Q
M1000 VPWR a_1226_296# a_1144_508# VPB pshort w=420000u l=180000u
+  ad=2.2454e+12p pd=1.922e+07u as=1.869e+11p ps=1.73e+06u
M1001 Q a_1226_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1002 VGND a_1226_296# Q VNB nlowvt w=740000u l=150000u
+  ad=1.88282e+12p pd=1.54e+07u as=4.44e+11p ps=4.16e+06u
M1003 Q a_1226_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_1226_296# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_654_503# a_27_74# a_547_485# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=1.6485e+11p ps=1.73e+06u
M1006 a_1144_508# a_209_368# a_1037_424# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.667e+11p ps=2.39e+06u
M1007 Q a_1226_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Q a_1226_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_440_503# D VPWR VPB pshort w=420000u l=180000u
+  ad=1.6485e+11p pd=1.73e+06u as=0p ps=0u
M1010 VPWR a_1226_296# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_696_458# a_547_485# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.98e+11p pd=1.97e+06u as=0p ps=0u
M1012 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1013 a_209_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1014 a_547_485# a_209_368# a_440_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1226_296# a_1037_424# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1016 VGND a_696_458# a_735_102# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 VGND a_1226_296# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1037_424# a_27_74# a_696_458# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.2e+11p ps=2.68e+06u
M1019 VPWR a_1037_424# a_1226_296# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1226_296# a_1178_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.323e+11p ps=1.47e+06u
M1021 a_735_102# a_209_368# a_547_485# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.51375e+11p ps=1.66e+06u
M1022 a_440_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1023 a_547_485# a_27_74# a_440_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1037_424# a_209_368# a_696_458# VNB nlowvt w=550000u l=150000u
+  ad=2.152e+11p pd=1.97e+06u as=0p ps=0u
M1025 a_209_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1026 VGND a_1037_424# a_1226_296# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1027 VPWR a_696_458# a_654_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1029 a_696_458# a_547_485# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1178_124# a_27_74# a_1037_424# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE ndiode p=7.32e+06u a=6.417e+11p
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
M1000 a_261_392# GATE VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=1.77765e+12p ps=1.19e+07u
M1001 a_477_124# a_309_338# a_83_260# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.692e+11p ps=2.3e+06u
M1002 VGND CLK a_315_54# VNB nlowvt w=740000u l=150000u
+  ad=1.19302e+12p pd=9.54e+06u as=2.183e+11p ps=2.07e+06u
M1003 a_83_260# a_309_338# a_261_392# VPB pshort w=1e+06u l=180000u
+  ad=3.676e+11p pd=3.06e+06u as=0p ps=0u
M1004 a_309_338# a_315_54# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 GCLK a_990_393# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1006 VPWR a_83_260# a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1007 a_487_508# a_315_54# a_83_260# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1008 VPWR CLK a_315_54# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 a_990_393# a_27_74# a_984_125# VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.536e+11p ps=1.76e+06u
M1010 VPWR a_27_74# a_487_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_27_74# a_990_393# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1012 a_984_125# CLK VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 GCLK a_990_393# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_309_338# a_315_54# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1015 a_990_393# CLK VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_27_74# a_477_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_83_260# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 a_267_80# GATE VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_83_260# a_315_54# a_267_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
M1000 a_83_244# a_315_338# a_267_392# VPB pshort w=1e+06u l=180000u
+  ad=4.054e+11p pd=3.24e+06u as=2.4e+11p ps=2.48e+06u
M1001 a_1044_387# CLK VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=2.5157e+12p ps=1.567e+07u
M1002 a_511_508# a_315_48# a_83_244# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1003 GCLK a_1044_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.45355e+12p ps=1.19e+07u
M1004 VPWR a_83_244# a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1005 VPWR a_27_74# a_1044_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_74# a_511_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_494_118# a_315_338# a_83_244# VNB nlowvt w=420000u l=150000u
+  ad=1.54875e+11p pd=1.7e+06u as=3.049e+11p ps=2.47e+06u
M1008 a_315_338# a_315_48# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1009 VGND a_1044_387# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_27_74# a_494_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_315_338# a_315_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 VPWR CLK a_315_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1013 a_83_244# a_315_48# a_267_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1014 a_267_74# GATE VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND CLK a_315_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 GCLK a_1044_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1017 a_1044_387# a_27_74# a_1044_119# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.554e+11p ps=1.9e+06u
M1018 VPWR a_1044_387# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1044_119# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_267_392# GATE VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_83_244# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
M1000 a_84_48# a_334_338# a_286_392# VPB pshort w=1e+06u l=180000u
+  ad=3.991e+11p pd=3.21e+06u as=2.4e+11p ps=2.48e+06u
M1001 VGND a_27_74# a_491_124# VNB nlowvt w=420000u l=150000u
+  ad=1.78525e+12p pd=1.468e+07u as=2.3775e+11p ps=2.39e+06u
M1002 VPWR a_27_74# a_527_508# VPB pshort w=420000u l=180000u
+  ad=3.0253e+12p pd=1.906e+07u as=1.008e+11p ps=1.32e+06u
M1003 VPWR a_84_48# a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1004 GCLK a_1047_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.216e+11p pd=5.59e+06u as=0p ps=0u
M1005 a_1047_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1006 GCLK a_1047_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 GCLK a_1047_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1047_368# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.416e+11p pd=2.85e+06u as=0p ps=0u
M1009 VGND a_1047_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_1047_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_491_124# a_334_338# a_84_48# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.587e+11p ps=2.25e+06u
M1012 VPWR CLK a_334_54# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 VGND a_1047_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_27_74# a_1047_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_334_338# a_334_54# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 GCLK a_1047_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_286_80# GATE VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1018 a_84_48# a_334_54# a_286_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND CLK a_334_54# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.333e+11p ps=2.19e+06u
M1020 VGND a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1021 a_1047_368# a_27_74# a_1047_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 VPWR a_1047_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_286_392# GATE VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_527_508# a_334_54# a_84_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_334_338# a_334_54# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.675e+11p pd=2.66e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR RESET_B a_889_92# VPB pshort w=1.12e+06u l=180000u
+  ad=2.18775e+12p pd=1.595e+07u as=3.136e+11p ps=2.8e+06u
M1001 a_608_74# a_27_424# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.4043e+12p ps=1.104e+07u
M1002 a_686_74# a_231_74# a_608_74# VNB nlowvt w=640000u l=150000u
+  ad=3.835e+11p pd=2.53e+06u as=0p ps=0u
M1003 a_231_74# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 a_805_508# a_231_74# a_686_74# VPB pshort w=420000u l=180000u
+  ad=2.121e+11p pd=1.85e+06u as=3.115e+11p ps=2.71e+06u
M1005 VGND RESET_B a_1133_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1006 a_686_74# a_373_74# a_614_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1007 a_231_74# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 VGND D a_27_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 Q_N a_1437_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1010 VGND a_889_92# a_1437_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.925e+11p ps=1.8e+06u
M1011 VPWR a_889_92# a_805_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR D a_27_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 a_889_92# a_686_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_841_118# a_373_74# a_686_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1015 VGND a_231_74# a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 Q a_889_92# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1017 a_1133_74# a_686_74# a_889_92# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 Q a_889_92# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 a_614_392# a_27_424# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q_N a_1437_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 VPWR a_889_92# a_1437_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1022 VPWR a_231_74# a_373_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=3.704e+11p ps=2.85e+06u
M1023 VGND a_889_92# a_841_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_838_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=2.6628e+12p pd=2.07e+07u as=3.024e+11p ps=2.78e+06u
M1001 a_1066_74# a_670_74# a_838_48# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.109e+11p ps=2.05e+06u
M1002 VGND RESET_B a_1066_74# VNB nlowvt w=740000u l=150000u
+  ad=1.80345e+12p pd=1.499e+07u as=0p ps=0u
M1003 Q a_838_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 VPWR a_838_48# a_786_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.869e+11p ps=1.73e+06u
M1005 VPWR a_230_74# a_363_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=3.704e+11p ps=2.85e+06u
M1006 a_592_74# a_27_112# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1007 a_670_74# a_230_74# a_592_74# VNB nlowvt w=640000u l=150000u
+  ad=2.44e+11p pd=2.18e+06u as=0p ps=0u
M1008 Q_N a_1448_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 a_598_392# a_27_112# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1010 VPWR a_1448_74# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_838_48# a_670_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1012 VPWR D a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 a_230_74# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_786_508# a_230_74# a_670_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.265e+11p ps=2.74e+06u
M1015 a_230_74# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 VGND D a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1017 a_790_74# a_363_74# a_670_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_1448_74# a_838_48# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1019 VGND a_838_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1448_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1021 a_1448_74# a_838_48# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1022 VGND a_230_74# a_363_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 VGND a_838_48# a_790_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_670_74# a_363_74# a_598_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_838_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR RESET_B a_838_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_1448_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 Q a_823_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.30975e+12p ps=1.109e+07u
M1001 a_643_80# a_226_104# a_567_392# VPB pshort w=1e+06u l=180000u
+  ad=3.315e+11p pd=2.75e+06u as=2.1e+11p ps=2.42e+06u
M1002 VGND D a_27_142# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1003 VGND a_226_104# a_353_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.59e+11p ps=2.18e+06u
M1004 VPWR a_823_98# a_1342_74# VPB pshort w=840000u l=180000u
+  ad=1.9237e+12p pd=1.499e+07u as=2.352e+11p ps=2.24e+06u
M1005 VPWR a_823_98# a_756_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1006 VGND a_823_98# a_775_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_571_80# a_27_142# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1008 a_643_80# a_353_98# a_571_80# VNB nlowvt w=640000u l=150000u
+  ad=2.692e+11p pd=2.3e+06u as=0p ps=0u
M1009 a_823_98# a_643_80# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1010 VGND a_823_98# a_1342_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1011 VPWR a_226_104# a_353_98# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1012 a_226_104# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.94e+11p pd=2.38e+06u as=0p ps=0u
M1013 VPWR RESET_B a_823_98# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q a_823_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 a_775_124# a_226_104# a_643_80# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_226_104# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.701e+11p pd=2.21e+06u as=0p ps=0u
M1017 VGND RESET_B a_1051_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1018 Q_N a_1342_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1019 a_756_508# a_353_98# a_643_80# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1051_74# a_643_80# a_823_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1021 a_567_392# a_27_142# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q_N a_1342_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.738e+11p pd=2.22e+06u as=0p ps=0u
M1023 VPWR D a_27_142# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR D a_27_112# VPB pshort w=840000u l=180000u
+  ad=2.6463e+12p pd=2.068e+07u as=2.352e+11p ps=2.24e+06u
M1001 VPWR a_230_74# a_363_82# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1002 VGND a_230_74# a_363_82# VNB nlowvt w=740000u l=150000u
+  ad=1.8561e+12p pd=1.54e+07u as=2.109e+11p ps=2.05e+06u
M1003 a_773_124# a_230_74# a_641_80# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.692e+11p ps=2.3e+06u
M1004 a_569_80# a_27_112# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1005 Q_N a_1449_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 VGND a_821_98# a_1449_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1007 VPWR a_821_98# a_760_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1008 VPWR a_1449_368# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND RESET_B a_1049_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1010 a_569_392# a_27_112# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1011 Q_N a_1449_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 VPWR a_821_98# a_1449_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1013 a_230_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_641_80# a_230_74# a_569_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=0p ps=0u
M1015 VGND D a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1016 a_1049_74# a_641_80# a_821_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_230_74# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.772e+11p pd=2.34e+06u as=0p ps=0u
M1018 VGND a_821_98# a_773_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_1449_368# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_760_508# a_363_82# a_641_80# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q a_821_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1022 VPWR a_821_98# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_641_80# a_363_82# a_569_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q a_821_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1025 VGND a_821_98# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR RESET_B a_821_98# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=2.88e+06u
M1027 a_821_98# a_641_80# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=1.64835e+12p ps=1.063e+07u
M1001 VGND a_897_406# a_854_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1002 Q a_897_406# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.70685e+12p ps=1.247e+07u
M1003 a_854_74# a_357_392# a_657_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.915e+11p ps=1.93e+06u
M1004 a_573_392# a_27_136# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1005 a_232_98# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1006 a_796_508# a_232_98# a_657_392# VPB pshort w=420000u l=180000u
+  ad=2.121e+11p pd=1.85e+06u as=3.816e+11p ps=3.03e+06u
M1007 VPWR a_897_406# a_796_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND RESET_B a_1139_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1009 VPWR a_232_98# a_357_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1010 a_681_74# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1011 VPWR RESET_B a_897_406# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.4e+11p ps=2.88e+06u
M1012 VPWR D a_27_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1014 a_1139_74# a_657_392# a_897_406# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1015 Q a_897_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.701e+11p pd=2.21e+06u as=0p ps=0u
M1016 VGND a_232_98# a_357_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_657_392# a_232_98# a_681_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_657_392# a_357_392# a_573_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_897_406# a_657_392# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 VGND RESET_B a_1153_74# VNB nlowvt w=740000u l=150000u
+  ad=2.30995e+12p pd=1.387e+07u as=1.776e+11p ps=1.96e+06u
M1001 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.257e+11p pd=2.09e+06u as=0p ps=0u
M1002 a_1153_74# a_673_392# a_913_406# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1003 a_589_392# a_27_136# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.6589e+12p ps=1.646e+07u
M1004 Q a_913_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VPWR a_913_406# a_781_504# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.772e+11p ps=2.16e+06u
M1006 Q a_913_406# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1007 VGND a_232_98# a_373_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1008 a_913_406# a_673_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1009 VPWR a_913_406# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_673_392# a_373_82# a_589_392# VPB pshort w=1e+06u l=180000u
+  ad=3.158e+11p pd=2.72e+06u as=0p ps=0u
M1011 a_232_98# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1012 a_781_504# a_232_98# a_673_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_913_406# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_673_392# a_232_98# a_697_74# VNB nlowvt w=640000u l=150000u
+  ad=1.915e+11p pd=1.93e+06u as=1.536e+11p ps=1.76e+06u
M1015 VPWR D a_27_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1016 a_697_74# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1018 VGND a_913_406# a_870_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1019 VPWR RESET_B a_913_406# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_870_74# a_373_82# a_673_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_232_98# a_373_82# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_750_504# a_232_98# a_642_392# VPB pshort w=420000u l=180000u
+  ad=2.898e+11p pd=2.22e+06u as=3.158e+11p ps=2.72e+06u
M1001 VGND a_888_406# Q VNB nlowvt w=740000u l=150000u
+  ad=2.1144e+12p pd=1.632e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_1035_74# RESET_B VGND VNB nlowvt w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=0p ps=0u
M1003 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1004 VGND a_888_406# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_564_392# a_27_136# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=2.5597e+12p ps=1.989e+07u
M1006 a_839_74# a_348_392# a_642_392# VNB nlowvt w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=1.915e+11p ps=1.93e+06u
M1007 a_232_98# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 VPWR a_232_98# a_348_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 a_1035_74# a_642_392# a_888_406# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1010 VPWR a_888_406# a_750_504# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_888_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_888_406# a_642_392# VPWR VPB pshort w=840000u l=180000u
+  ad=5.124e+11p pd=4.58e+06u as=0p ps=0u
M1013 VPWR D a_27_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1014 a_888_406# RESET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_888_406# a_839_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_642_392# a_888_406# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_642_392# a_232_98# a_666_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1018 a_666_74# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_888_406# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=7.168e+11p ps=5.76e+06u
M1020 VGND a_232_98# a_348_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1021 VGND RESET_B a_1035_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q a_888_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_888_406# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1025 Q a_888_406# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_888_406# a_642_392# a_1035_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_888_406# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_642_392# a_348_392# a_564_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR RESET_B a_888_406# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_643_74# a_219_424# a_571_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR a_219_424# a_363_74# VPB pshort w=840000u l=180000u
+  ad=1.4754e+12p pd=1.132e+07u as=2.352e+11p ps=2.24e+06u
M1002 VPWR RESET_B a_817_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1003 a_817_48# a_643_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Q a_817_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 a_762_508# a_363_74# a_643_74# VPB pshort w=420000u l=180000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1006 a_219_424# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=4.2675e+11p pd=2.84e+06u as=0p ps=0u
M1007 a_219_424# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=9.349e+11p ps=8.16e+06u
M1008 VPWR D a_27_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 VGND RESET_B a_1045_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1010 a_769_74# a_219_424# a_643_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.907e+11p ps=2.24e+06u
M1011 VGND a_817_48# a_769_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_219_424# a_363_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.2225e+11p ps=2.64e+06u
M1013 VPWR a_817_48# a_762_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q a_817_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1015 a_1045_74# a_643_74# a_817_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 a_571_392# a_27_424# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND D a_27_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1018 a_565_74# a_27_424# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_643_74# a_363_74# a_565_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_759_508# a_347_98# a_646_74# VPB pshort w=420000u l=180000u
+  ad=2.121e+11p pd=1.85e+06u as=3.115e+11p ps=2.71e+06u
M1001 VGND a_235_74# a_347_98# VNB nlowvt w=740000u l=150000u
+  ad=1.38725e+12p pd=1.126e+07u as=2.701e+11p ps=2.21e+06u
M1002 VPWR D a_27_392# VPB pshort w=840000u l=180000u
+  ad=2.11845e+12p pd=1.561e+07u as=2.352e+11p ps=2.24e+06u
M1003 a_568_74# a_27_392# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1004 a_646_74# a_347_98# a_568_74# VNB nlowvt w=640000u l=150000u
+  ad=3.21575e+11p pd=2.36e+06u as=0p ps=0u
M1005 VGND RESET_B a_1060_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1006 Q a_832_55# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=0p ps=0u
M1007 VPWR a_235_74# a_347_98# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1008 Q a_832_55# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1009 a_832_55# a_646_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1010 VPWR RESET_B a_832_55# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_832_55# a_759_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_27_392# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 VPWR a_832_55# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_568_392# a_27_392# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1015 a_235_74# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 a_646_74# a_235_74# a_568_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1060_74# a_646_74# a_832_55# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 VGND a_832_55# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_784_81# a_235_74# a_646_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1020 VGND a_832_55# a_784_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_235_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 VPWR D a_27_126# VPB pshort w=840000u l=180000u
+  ad=2.5342e+12p pd=2.013e+07u as=2.352e+11p ps=2.24e+06u
M1001 a_938_74# a_640_74# a_797_48# VNB nlowvt w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=1.824e+11p ps=1.85e+06u
M1002 a_559_74# a_27_126# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.632e+11p pd=1.79e+06u as=1.6158e+12p ps=1.463e+07u
M1003 a_755_74# a_243_394# a_640_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.555e+11p ps=2.13e+06u
M1004 VPWR a_797_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.832e+11p ps=5.7e+06u
M1005 a_243_394# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 VPWR a_243_394# a_364_120# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1007 a_797_48# a_640_74# a_938_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_797_48# a_640_74# VPWR VPB pshort w=840000u l=180000u
+  ad=4.956e+11p pd=4.54e+06u as=0p ps=0u
M1009 Q a_797_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1010 Q a_797_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR RESET_B a_797_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_640_74# a_797_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_797_48# RESET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_797_48# a_750_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.869e+11p ps=1.73e+06u
M1015 a_640_74# a_243_394# a_565_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=2.1e+11p ps=2.42e+06u
M1016 a_243_394# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.814e+11p pd=2.35e+06u as=0p ps=0u
M1017 VGND D a_27_126# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1018 VGND RESET_B a_938_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Q a_797_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_797_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_243_394# a_364_120# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1022 Q a_797_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_797_48# a_755_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_797_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_750_508# a_364_120# a_640_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_640_74# a_364_120# a_559_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_565_392# a_27_126# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_938_74# RESET_B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_797_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
M1000 VPWR D a_27_120# VPB pshort w=840000u l=180000u
+  ad=1.6835e+12p pd=1.404e+07u as=2.814e+11p ps=2.35e+06u
M1001 a_232_82# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1002 a_574_392# a_27_120# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1003 a_232_82# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.4754e+12p ps=1.217e+07u
M1004 VGND a_863_294# a_852_123# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 a_863_294# a_653_79# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.183e+11p pd=2.07e+06u as=0p ps=0u
M1006 a_808_392# a_232_82# a_653_79# VPB pshort w=420000u l=180000u
+  ad=1.281e+11p pd=1.45e+06u as=3.844e+11p ps=3.14e+06u
M1007 Q_N a_1350_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 VGND a_232_82# a_343_80# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.182e+11p ps=2.34e+06u
M1009 VGND a_863_294# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1010 a_852_123# a_343_80# a_653_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.099e+11p ps=2.97e+06u
M1011 VPWR a_863_294# a_808_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_653_79# a_232_82# a_575_79# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1013 a_575_79# a_27_120# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_653_79# a_343_80# a_574_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_863_294# a_653_79# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1016 a_1350_424# a_863_294# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1017 a_1350_424# a_863_294# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1018 Q_N a_1350_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1019 VPWR a_863_294# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1020 VGND D a_27_120# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1021 VPWR a_232_82# a_343_80# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_887_270# Q VPB pshort w=1.12e+06u l=180000u
+  ad=2.3791e+12p pd=1.953e+07u as=3.024e+11p ps=2.78e+06u
M1001 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.0325e+12p ps=1.669e+07u
M1002 Q a_887_270# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 Q_N a_1442_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1004 VGND a_232_98# a_343_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.817e+11p ps=2.29e+06u
M1005 VPWR a_1442_94# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_817_392# a_232_98# a_647_79# VPB pshort w=420000u l=180000u
+  ad=1.47e+11p pd=1.54e+06u as=4.159e+11p ps=3.29e+06u
M1007 Q_N a_1442_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 VGND a_887_270# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_887_270# a_647_79# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1010 a_1442_94# a_887_270# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1011 a_568_392# a_27_136# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1012 a_569_79# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1013 a_647_79# a_232_98# a_569_79# VNB nlowvt w=640000u l=150000u
+  ad=3.952e+11p pd=2.9e+06u as=0p ps=0u
M1014 VGND a_1442_94# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_887_270# a_647_79# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 a_1442_94# a_887_270# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1017 a_647_79# a_343_74# a_568_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1019 a_232_98# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1020 VPWR D a_27_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=3.066e+11p ps=2.41e+06u
M1021 VPWR a_887_270# a_817_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_887_270# a_839_123# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1023 VPWR a_232_98# a_343_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1024 Q a_887_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_839_123# a_343_74# a_647_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_231_74# a_373_82# VPB pshort w=840000u l=180000u
+  ad=1.95315e+12p pd=1.524e+07u as=2.352e+11p ps=2.24e+06u
M1001 a_589_392# a_27_413# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1002 a_231_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.4685e+12p ps=1.184e+07u
M1003 a_815_124# a_231_74# a_667_80# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.028e+11p ps=2.46e+06u
M1004 a_863_98# a_667_80# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 VGND D a_27_413# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1006 VPWR a_863_98# a_773_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1007 a_863_98# a_667_80# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 Q_N a_1350_116# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 Q_N a_1350_116# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1010 VPWR D a_27_413# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1011 a_667_80# a_373_82# a_589_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1012 a_589_80# a_27_413# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_231_74# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1014 a_1350_116# a_863_98# VPWR VPB pshort w=840000u l=180000u
+  ad=2.31e+11p pd=2.23e+06u as=0p ps=0u
M1015 VGND a_863_98# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1016 a_667_80# a_231_74# a_589_392# VPB pshort w=1e+06u l=180000u
+  ad=3.065e+11p pd=2.7e+06u as=0p ps=0u
M1017 VPWR a_863_98# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1018 a_1350_116# a_863_98# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1019 VGND a_231_74# a_373_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1020 VGND a_863_98# a_815_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_773_508# a_373_82# a_667_80# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
M1000 a_815_508# a_220_419# a_672_392# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=4.915e+11p ps=3.07e+06u
M1001 Q a_863_441# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=1.31878e+12p ps=1.016e+07u
M1002 Q a_863_441# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.48785e+12p ps=1.153e+07u
M1003 VGND a_220_419# a_369_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 a_588_392# a_27_115# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1005 VGND D a_27_115# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1006 a_863_441# a_672_392# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1007 a_871_139# a_369_392# a_672_392# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.786e+11p ps=2.52e+06u
M1008 a_672_392# a_369_392# a_588_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_220_419# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 VPWR a_863_441# a_815_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_220_419# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=3.066e+11p pd=2.41e+06u as=0p ps=0u
M1012 VGND a_863_441# a_871_139# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_863_441# a_672_392# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1014 VPWR D a_27_115# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1015 VPWR a_220_419# a_369_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1016 a_655_79# a_27_115# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1017 a_672_392# a_220_419# a_655_79# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
M1000 Q a_842_405# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=1.54015e+12p ps=1.207e+07u
M1001 VPWR D a_27_120# VPB pshort w=840000u l=180000u
+  ad=1.89385e+12p pd=1.485e+07u as=2.352e+11p ps=2.24e+06u
M1002 a_672_392# a_232_82# a_658_79# VNB nlowvt w=640000u l=150000u
+  ad=2.803e+11p pd=2.53e+06u as=1.536e+11p ps=1.76e+06u
M1003 a_658_79# a_27_120# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_232_82# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VPWR a_842_405# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.528e+11p ps=2.87e+06u
M1006 VGND a_842_405# a_875_139# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 VPWR a_842_405# a_794_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VGND a_232_82# a_369_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_588_392# a_27_120# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1010 VGND a_842_405# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_842_405# a_672_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_672_392# a_369_392# a_588_392# VPB pshort w=1e+06u l=180000u
+  ad=3.83875e+11p pd=2.86e+06u as=0p ps=0u
M1013 a_875_139# a_369_392# a_672_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_842_405# a_672_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 a_794_503# a_232_82# a_672_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND D a_27_120# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1017 a_232_82# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1018 VPWR a_232_82# a_369_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1019 Q a_842_405# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
M1000 a_792_508# a_232_114# a_678_392# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=3.262e+11p ps=2.78e+06u
M1001 a_678_392# a_232_114# a_658_79# VNB nlowvt w=640000u l=150000u
+  ad=3.259e+11p pd=2.57e+06u as=1.536e+11p ps=1.76e+06u
M1002 a_658_79# a_27_115# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.78397e+12p ps=1.439e+07u
M1003 VGND a_840_395# a_895_123# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 a_840_395# a_678_392# VPWR VPB pshort w=840000u l=180000u
+  ad=2.73e+11p pd=2.33e+06u as=2.1628e+12p ps=1.704e+07u
M1005 VGND a_232_114# a_369_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1006 a_232_114# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1007 VGND a_678_392# a_840_395# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1008 a_895_123# a_369_392# a_678_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_678_392# a_369_392# a_594_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1010 VGND D a_27_115# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1011 VPWR D a_27_115# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1012 Q a_840_395# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.888e+11p pd=5.71e+06u as=0p ps=0u
M1013 Q a_840_395# VGND VNB nlowvt w=740000u l=150000u
+  ad=5.143e+11p pd=4.35e+06u as=0p ps=0u
M1014 VPWR a_840_395# a_792_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_840_395# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_232_114# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1017 VPWR a_840_395# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_840_395# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_840_395# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_232_114# a_369_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1021 a_594_392# a_27_115# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_678_392# a_840_395# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_840_395# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_840_395# a_678_392# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_840_395# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxtp_1 D GATE VGND VNB VPB VPWR Q
M1000 Q a_386_326# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.60698e+12p ps=1.245e+07u
M1001 VGND a_119_88# a_239_85# VNB nlowvt w=740000u l=150000u
+  ad=1.47895e+12p pd=1.06e+07u as=4.458e+11p ps=4.22e+06u
M1002 a_422_392# a_386_326# VPWR VPB pshort w=420000u l=180000u
+  ad=3.0425e+11p pd=3.2e+06u as=0p ps=0u
M1003 a_685_59# a_562_123# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 a_592_149# a_562_123# a_514_149# VNB nlowvt w=420000u l=150000u
+  ad=2.753e+11p pd=2.41e+06u as=1.008e+11p ps=1.32e+06u
M1005 Q a_386_326# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 a_119_88# D VGND VNB nlowvt w=550000u l=150000u
+  ad=1.815e+11p pd=1.76e+06u as=0p ps=0u
M1007 VPWR a_119_88# a_229_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1008 a_119_88# D VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1009 VGND a_592_149# a_386_326# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1010 VPWR a_592_149# a_386_326# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.528e+11p ps=2.87e+06u
M1011 a_685_59# a_562_123# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1012 VPWR GATE a_562_123# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 a_592_149# a_562_123# a_229_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=0p ps=0u
M1014 a_514_149# a_386_326# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_239_85# a_685_59# a_592_149# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND GATE a_562_123# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.22e+11p ps=2.08e+06u
M1017 a_422_392# a_685_59# a_592_149# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlygate4sd1_1 A VGND VNB VPB VPWR X
M1000 VPWR a_288_74# a_405_138# VPB pshort w=1e+06u l=180000u
+  ad=9.874e+11p pd=6.28e+06u as=5.8e+11p ps=3.16e+06u
M1001 X a_405_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1002 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1003 VGND a_288_74# a_405_138# VNB nlowvt w=420000u l=150000u
+  ad=5.384e+11p pd=4.48e+06u as=2.562e+11p ps=2.06e+06u
M1004 VPWR A a_28_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 X a_405_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1007 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlygate4sd2_1 A VGND VNB VPB VPWR X
M1000 X a_405_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=9.174e+11p ps=6.14e+06u
M1001 VPWR A a_28_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=5.258e+11p ps=4.42e+06u
M1003 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VGND a_288_74# a_405_138# VNB nlowvt w=420000u l=180000u
+  ad=0p pd=0u as=2.436e+11p ps=2e+06u
M1005 X a_405_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1006 VPWR a_288_74# a_405_138# VPB pshort w=1e+06u l=250000u
+  ad=0p pd=0u as=5.1e+11p ps=3.02e+06u
M1007 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=250000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlygate4sd3_1 A VGND VNB VPB VPWR X
M1000 X a_405_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=6.674e+11p ps=5.64e+06u
M1001 a_289_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=5.279e+11p ps=4.43e+06u
M1002 VPWR a_289_74# a_405_138# VPB pshort w=1e+06u l=500000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1003 a_289_74# a_28_74# VPWR VPB pshort w=1e+06u l=500000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1004 VPWR A a_28_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 VGND a_289_74# a_405_138# VNB nlowvt w=420000u l=180000u
+  ad=0p pd=0u as=2.436e+11p ps=2e+06u
M1007 X a_405_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlymetal6s2s_1 A VGND VNB VPB VPWR X
M1000 VPWR A a_28_138# VPB pshort w=420000u l=180000u
+  ad=9.737e+11p pd=8.74e+06u as=1.092e+11p ps=1.36e+06u
M1001 VGND a_497_74# a_604_138# VNB nlowvt w=420000u l=150000u
+  ad=6.828e+11p pd=6.48e+06u as=1.113e+11p ps=1.37e+06u
M1002 X a_28_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1003 X a_28_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1004 VPWR X a_316_138# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 a_785_74# a_604_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1006 VGND A a_28_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VGND X a_316_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_497_74# a_316_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1009 a_497_74# a_316_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1010 VPWR a_497_74# a_604_138# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 a_785_74# a_604_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlymetal6s4s_1 A VGND VNB VPB VPWR X
M1000 VPWR A a_28_138# VPB pshort w=420000u l=180000u
+  ad=9.737e+11p pd=8.74e+06u as=1.092e+11p ps=1.36e+06u
M1001 VGND X a_604_138# VNB nlowvt w=420000u l=150000u
+  ad=6.828e+11p pd=6.48e+06u as=1.113e+11p ps=1.37e+06u
M1002 a_209_74# a_28_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1003 a_209_74# a_28_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1004 VPWR a_209_74# a_316_138# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 a_785_74# a_604_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1006 VGND A a_28_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VGND a_209_74# a_316_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 X a_316_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1009 X a_316_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1010 VPWR X a_604_138# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 a_785_74# a_604_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlymetal6s6s_1 A VGND VNB VPB VPWR X
M1000 VPWR A a_28_138# VPB pshort w=420000u l=180000u
+  ad=9.737e+11p pd=8.74e+06u as=1.092e+11p ps=1.36e+06u
M1001 VGND a_497_74# a_604_138# VNB nlowvt w=420000u l=150000u
+  ad=6.828e+11p pd=6.48e+06u as=1.113e+11p ps=1.37e+06u
M1002 a_209_74# a_28_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1003 a_209_74# a_28_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1004 VPWR a_209_74# a_316_138# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 X a_604_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1006 VGND A a_28_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VGND a_209_74# a_316_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_497_74# a_316_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1009 a_497_74# a_316_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1010 VPWR a_497_74# a_604_138# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 X a_604_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ebufn_1 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_27_404# VPB pshort w=840000u l=180000u
+  ad=7.441e+11p pd=5.78e+06u as=2.352e+11p ps=2.24e+06u
M1001 a_569_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1002 a_229_74# A VGND VNB nlowvt w=550000u l=150000u
+  ad=1.4575e+11p pd=1.63e+06u as=3.759e+11p ps=3.75e+06u
M1003 a_229_74# A VPWR VPB pshort w=840000u l=180000u
+  ad=2.436e+11p pd=2.26e+06u as=0p ps=0u
M1004 Z a_229_74# a_569_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 a_569_74# a_27_404# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1006 Z a_229_74# a_569_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VGND TE_B a_27_404# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ebufn_2 A TE_B VGND VNB VPB VPWR Z
M1000 a_84_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=4.797e+11p ps=4.17e+06u
M1001 VPWR TE_B a_283_48# VPB pshort w=1e+06u l=180000u
+  ad=1.0179e+12p pd=6.44e+06u as=2.8e+11p ps=2.56e+06u
M1002 VGND a_283_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=7.289e+11p ps=6.41e+06u
M1003 a_27_74# a_283_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR TE_B a_33_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=9.856e+11p ps=8.48e+06u
M1005 a_33_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=2.88e+06u
M1006 a_33_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z a_84_48# a_33_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1009 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_84_48# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1011 VGND TE_B a_283_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ebufn_4 A TE_B VGND VNB VPB VPWR Z
M1000 Z a_27_368# a_348_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.5288e+12p ps=1.393e+07u
M1001 a_208_74# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=9.352e+11p ps=8.39e+06u
M1002 a_348_368# a_27_368# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Z a_27_368# a_348_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=2.109e+11p ps=2.05e+06u
M1005 a_378_74# a_27_368# Z VNB nlowvt w=740000u l=150000u
+  ad=1.0323e+12p pd=1.019e+07u as=4.292e+11p ps=4.12e+06u
M1006 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1007 VGND a_208_74# a_378_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_378_74# a_208_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_208_74# a_378_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_348_368# a_27_368# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_208_74# TE_B VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_378_74# a_27_368# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR TE_B a_348_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Z a_27_368# a_378_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_378_74# a_208_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_348_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR TE_B a_348_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Z a_27_368# a_378_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_348_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ebufn_8 A TE_B VGND VNB VPB VPWR Z
M1000 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.0054e+12p pd=1.874e+07u as=1.2506e+12p ps=1.226e+07u
M1001 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.3048e+12p pd=1.129e+07u as=2.8168e+12p ps=2.519e+07u
M1002 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=9.213e+11p ps=8.41e+06u
M1008 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.4573e+12p ps=1.808e+07u
M1010 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_84_48# A VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A a_84_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_84_48# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR TE_B a_833_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.544e+11p ps=3.23e+06u
M1029 VGND TE_B a_833_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1030 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR A a_84_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
M1000 a_1198_97# a_1008_74# a_27_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.349e+11p ps=4.69e+06u
M1001 a_527_74# a_161_446# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.908e+12p ps=1.641e+07u
M1002 a_27_74# a_575_48# a_527_74# VNB nlowvt w=420000u l=150000u
+  ad=4.158e+11p pd=4.5e+06u as=0p ps=0u
M1003 a_2209_443# a_1008_74# a_1879_74# VPB pshort w=420000u l=180000u
+  ad=1.26e+11p pd=1.44e+06u as=3.262e+11p ps=2.78e+06u
M1004 a_1807_74# a_1419_71# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1005 a_1419_71# a_1198_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=2.42065e+12p ps=2.12e+07u
M1006 a_1879_74# a_1008_74# a_1807_74# VNB nlowvt w=740000u l=150000u
+  ad=7.478e+11p pd=4.66e+06u as=0p ps=0u
M1007 a_1426_508# a_818_74# a_1198_97# VPB pshort w=420000u l=180000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1008 VPWR DE a_161_446# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1009 a_559_504# DE VPWR VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VGND a_575_48# a_2227_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1011 VPWR a_161_446# a_119_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 a_2011_392# a_1419_71# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1013 a_575_48# a_1879_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1014 a_1334_97# a_1008_74# a_1198_97# VNB nlowvt w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=2.226e+11p ps=1.9e+06u
M1015 a_1419_71# a_1198_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1016 a_575_48# a_1879_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1017 VGND a_1879_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 VGND DE a_145_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 VGND a_1419_71# a_1334_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q_N a_575_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_2227_118# a_818_74# a_1879_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_575_48# a_2209_443# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_1419_71# a_1426_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND DE a_161_446# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.281e+11p ps=1.45e+06u
M1025 a_818_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1026 VPWR a_1879_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1027 a_119_508# D a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1008_74# a_818_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1029 a_1008_74# a_818_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1030 Q_N a_575_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1031 a_818_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1032 a_145_74# D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_74# a_575_48# a_559_504# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1198_97# a_818_74# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1879_74# a_818_74# a_2011_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
M1000 VPWR a_533_61# a_2091_502# VPB pshort w=420000u l=180000u
+  ad=2.10553e+12p pd=1.949e+07u as=1.008e+11p ps=1.32e+06u
M1001 VGND a_1409_64# a_1349_90# VNB nlowvt w=420000u l=150000u
+  ad=1.8056e+12p pd=1.622e+07u as=1.26e+11p ps=1.44e+06u
M1002 VGND a_533_61# a_1997_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1003 a_533_61# a_1895_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1004 a_1409_64# a_1156_90# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1005 a_958_74# a_763_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1006 VGND DE a_131_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_1997_74# a_763_74# a_1895_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.424e+11p ps=2.2e+06u
M1008 a_117_508# D a_27_508# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=3.339e+11p ps=4.11e+06u
M1009 a_131_74# D a_27_508# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.591e+11p ps=4.23e+06u
M1010 VGND DE a_159_446# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1011 a_763_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=0p ps=0u
M1012 a_1797_74# a_1409_64# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1013 a_1156_90# a_958_74# a_27_508# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1014 a_533_61# a_1895_74# VPWR VPB pshort w=640000u l=180000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1015 VPWR a_159_446# a_117_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_557_436# DE VPWR VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1017 a_1385_508# a_763_74# a_1156_90# VPB pshort w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1018 a_1797_392# a_1409_64# VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.55e+11p pd=3.51e+06u as=0p ps=0u
M1019 VGND a_1895_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1020 VPWR a_1409_64# a_1385_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_491_87# a_159_446# VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1022 a_27_508# a_533_61# a_491_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1409_64# a_1156_90# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1024 a_1156_90# a_763_74# a_27_508# VNB nlowvt w=420000u l=150000u
+  ad=3.423e+11p pd=2.47e+06u as=0p ps=0u
M1025 a_763_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1026 a_2091_502# a_958_74# a_1895_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.115e+11p ps=2.71e+06u
M1027 a_27_508# a_533_61# a_557_436# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1349_90# a_958_74# a_1156_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1895_74# a_958_74# a_1797_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1895_74# a_763_74# a_1797_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_1895_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1032 VPWR DE a_159_446# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1033 a_958_74# a_763_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvn_1 A TE_B VGND VNB VPB VPWR Z
M1000 a_281_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=3.616e+11p ps=2.95e+06u
M1001 Z A a_281_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_281_100# a_22_46# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.564e+11p ps=2.36e+06u
M1003 Z A a_281_100# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 VPWR TE_B a_22_46# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1005 VGND TE_B a_22_46# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvn_2 A TE_B VGND VNB VPB VPWR Z
M1000 VGND a_117_74# a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=3.269e+11p pd=3.45e+06u as=6.176e+11p ps=6.17e+06u
M1001 a_231_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1002 VPWR TE_B a_227_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.784e+11p pd=4.61e+06u as=9.296e+11p ps=8.38e+06u
M1003 a_227_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Z A a_227_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 a_227_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_117_74# TE_B VPWR VPB pshort w=640000u l=180000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1007 a_231_74# a_117_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_74# TE_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvn_4 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.744e+11p pd=8.46e+06u as=1.5344e+12p ps=1.394e+07u
M1001 a_281_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=1.0508e+12p pd=1.024e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_241_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_281_74# a_114_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=6.253e+11p ps=6.13e+06u
M1004 VPWR TE_B a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_241_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_114_74# a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_281_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1009 a_241_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Z A a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_241_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Z A a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_281_74# a_114_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_114_74# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 a_114_74# TE_B VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 Z A a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_114_74# a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvn_8 A TE_B VGND VNB VPB VPWR Z
M1000 a_239_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=2.744e+12p pd=2.506e+07u as=1.2656e+12p ps=1.122e+07u
M1001 Z A a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_126_74# TE_B VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.1433e+12p ps=1.049e+07u
M1003 a_293_74# a_126_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.924e+12p pd=1.852e+07u as=0p ps=0u
M1004 Z A a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_126_74# a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Z A a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=9.324e+11p pd=8.44e+06u as=0p ps=0u
M1007 a_239_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_126_74# a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_126_74# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.8592e+12p ps=1.452e+07u
M1010 Z A a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Z A a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_239_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z A a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Z A a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_293_74# a_126_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_126_74# a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_239_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_293_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR TE_B a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_239_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_239_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_126_74# a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR TE_B a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_293_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR TE_B a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_239_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_293_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR TE_B a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_293_74# a_126_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_293_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_293_74# a_126_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Z A a_239_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_239_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvp_1 A TE VGND VNB VPB VPWR Z
M1000 a_313_392# a_44_549# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=3.115e+11p ps=2.71e+06u
M1001 a_318_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.276e+11p ps=2.16e+06u
M1002 Z A a_318_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 VGND TE a_44_549# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.604e+11p ps=2.08e+06u
M1004 Z A a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1005 VPWR TE a_44_549# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.583e+11p ps=2.07e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvp_2 A TE VGND VNB VPB VPWR Z
M1000 VGND TE a_263_323# VNB nlowvt w=420000u l=150000u
+  ad=3.332e+11p pd=3.48e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_36_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=2.072e+11p ps=2.04e+06u
M1002 VPWR TE a_263_323# VPB pshort w=640000u l=180000u
+  ad=4.816e+11p pd=4.62e+06u as=1.76e+11p ps=1.83e+06u
M1003 Z A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=9.24e+11p ps=8.37e+06u
M1004 a_27_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_263_323# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_368# a_263_323# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND TE a_36_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_36_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z A a_36_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvp_4 A TE VGND VNB VPB VPWR Z
M1000 Z A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.552e+11p pd=5.65e+06u as=1.652e+12p ps=1.415e+07u
M1001 VGND TE a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=8.843e+11p pd=6.83e+06u as=1.1655e+12p ps=1.055e+07u
M1002 Z A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_473_323# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.856e+11p pd=8.48e+06u as=0p ps=0u
M1005 a_27_368# a_473_323# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.995e+11p ps=4.31e+06u
M1008 VPWR a_473_323# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR TE a_473_323# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1013 Z A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND TE a_473_323# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1015 a_27_368# a_473_323# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Z A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND TE a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvp_8 A TE VGND VNB VPB VPWR Z
M1000 VPWR a_802_323# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.512e+12p pd=1.39e+07u as=2.7328e+12p ps=2.504e+07u
M1001 VGND TE a_802_323# VNB nlowvt w=740000u l=150000u
+  ad=1.1433e+12p pd=1.049e+07u as=2.146e+11p ps=2.06e+06u
M1002 a_27_368# a_802_323# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_802_323# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.0276e+12p pd=1.88e+07u as=0p ps=0u
M1005 a_27_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=9.842e+11p ps=8.58e+06u
M1006 Z A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.2096e+12p ps=1.112e+07u
M1010 a_27_368# a_802_323# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND TE a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Z A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_802_323# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Z A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Z A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_368# a_802_323# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Z A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_802_323# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Z A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_368# a_802_323# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR TE a_802_323# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1026 a_27_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Z A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Z A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_27_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND TE a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND TE a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND TE a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_315_75# B a_237_75# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_69_260# CIN a_315_75# VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1002 a_936_75# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.65875e+12p ps=1.244e+07u
M1003 a_321_389# B a_220_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6175e+11p pd=3.07e+06u as=3.43375e+11p ps=2.86e+06u
M1004 a_69_260# CIN a_321_389# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 VPWR CIN a_512_347# VPB pshort w=1e+06u l=180000u
+  ad=2.0852e+12p pd=1.495e+07u as=6.3e+11p ps=5.26e+06u
M1006 a_512_347# a_465_249# a_69_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 COUT a_465_249# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1008 VGND CIN a_501_75# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.096e+11p ps=3.84e+06u
M1009 a_1110_347# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.35e+11p pd=5.47e+06u as=0p ps=0u
M1010 a_501_75# a_465_249# a_69_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_237_75# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_512_347# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_465_249# B a_919_347# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=3.25e+11p ps=2.65e+06u
M1014 VGND B a_501_75# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1100_75# B VGND VNB nlowvt w=640000u l=150000u
+  ad=8.888e+11p pd=5.27e+06u as=0p ps=0u
M1016 a_501_75# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_465_249# B a_936_75# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1018 COUT a_465_249# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1019 a_919_347# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1110_347# CIN a_465_249# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_69_260# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1022 VPWR A a_1110_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A a_1100_75# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1100_75# CIN a_465_249# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B a_512_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_69_260# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1027 a_220_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 VPWR B a_686_347# VPB pshort w=1e+06u l=180000u
+  ad=2.63765e+12p pd=1.825e+07u as=6.22125e+11p ps=5.5e+06u
M1001 a_995_347# a_339_347# a_701_79# VNB nlowvt w=740000u l=150000u
+  ad=2.59e+11p pd=2.18e+06u as=5.18e+11p ps=4.36e+06u
M1002 a_1205_79# B a_1119_79# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.072e+11p ps=2.04e+06u
M1003 VGND A a_1205_79# VNB nlowvt w=740000u l=150000u
+  ad=2.36723e+12p pd=1.592e+07u as=0p ps=0u
M1004 COUT a_339_347# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 a_27_79# B VGND VNB nlowvt w=740000u l=150000u
+  ad=6.327e+11p pd=4.67e+06u as=0p ps=0u
M1006 SUM a_995_347# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1007 COUT a_339_347# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=4.088e+11p pd=2.97e+06u as=0p ps=0u
M1008 VPWR A a_1205_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1009 a_686_347# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_339_347# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 SUM a_995_347# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1012 VGND a_339_347# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_27_378# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.5e+11p ps=5.1e+06u
M1014 a_27_378# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_995_347# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_995_347# a_339_347# a_686_347# VPB pshort w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=0p ps=0u
M1017 VPWR a_995_347# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B a_701_79# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_339_347# CIN a_27_378# VPB pshort w=1e+06u l=180000u
+  ad=5.6e+11p pd=3.12e+06u as=0p ps=0u
M1020 a_1097_347# CIN a_995_347# VPB pshort w=1e+06u l=180000u
+  ad=3.747e+11p pd=2.93e+06u as=0p ps=0u
M1021 a_701_79# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_487_347# B a_339_347# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1023 VGND A a_27_79# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1119_79# CIN a_995_347# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A a_487_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_686_347# CIN VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A a_487_79# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1028 a_487_79# B a_339_347# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.59e+11p ps=2.18e+06u
M1029 a_1205_368# B a_1097_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_339_347# CIN a_27_79# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_701_79# CIN VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 VPWR a_418_74# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=2.97415e+12p pd=2.322e+07u as=6.048e+11p ps=5.56e+06u
M1001 a_418_74# CIN a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=4.181e+11p ps=4.09e+06u
M1002 VGND A a_1238_74# VNB nlowvt w=740000u l=150000u
+  ad=2.9966e+12p pd=2.115e+07u as=2.664e+11p ps=2.2e+06u
M1003 VPWR A a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.23132e+12p ps=6.6e+06u
M1004 a_740_347# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1005 VPWR A a_538_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1006 a_740_347# CIN VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 SUM a_1024_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1008 SUM a_1024_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1144_347# CIN a_1024_74# VPB pshort w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=3.2e+11p ps=2.64e+06u
M1010 VPWR a_1024_74# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 COUT a_418_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1012 VPWR B a_740_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1024_74# a_418_74# a_740_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_418_74# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_734_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1016 a_1024_74# a_418_74# a_734_74# VNB nlowvt w=740000u l=150000u
+  ad=3.922e+11p pd=2.54e+06u as=0p ps=0u
M1017 a_27_392# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_1238_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.747e+11p ps=2.93e+06u
M1019 COUT a_418_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1024_74# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 COUT a_418_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1024_74# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1023 VPWR a_418_74# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 SUM a_1024_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 COUT a_418_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_532_74# B a_418_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1027 a_418_74# CIN a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1028 a_1160_74# CIN a_1024_74# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1029 a_538_347# B a_418_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1238_347# B a_1144_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_734_74# CIN VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND B a_734_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND A a_532_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_1024_74# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_418_74# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 SUM a_1024_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1238_74# B a_1160_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_231_132# CI VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.06802e+12p pd=6.52e+06u as=2.27012e+12p ps=1.57e+07u
M1001 a_410_58# a_811_379# a_879_55# VNB nlowvt w=640000u l=150000u
+  ad=2.6395e+11p pd=2.41e+06u as=4.9405e+11p ps=5.22e+06u
M1002 a_83_21# a_811_379# a_231_132# VNB nlowvt w=640000u l=150000u
+  ad=2.375e+11p pd=2.16e+06u as=3.808e+11p ps=3.75e+06u
M1003 a_644_104# a_231_132# VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.31125e+11p pd=3.21e+06u as=0p ps=0u
M1004 a_811_379# a_879_55# a_1852_374# VNB nlowvt w=640000u l=150000u
+  ad=6.528e+11p pd=3.32e+06u as=5.128e+11p ps=4.25e+06u
M1005 a_1023_379# a_879_55# a_1852_374# VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=1.57615e+12p ps=7.29e+06u
M1006 a_1023_379# a_879_55# a_1660_374# VNB nlowvt w=640000u l=150000u
+  ad=4.965e+11p pd=2.98e+06u as=5.157e+11p ps=4.37e+06u
M1007 VPWR a_410_58# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.5085e+11p ps=3.26e+06u
M1008 VGND a_410_58# COUT VNB nlowvt w=740000u l=150000u
+  ad=1.8144e+12p pd=1.292e+07u as=2.072e+11p ps=2.04e+06u
M1009 a_1660_374# B a_1023_379# VPB pshort w=840000u l=180000u
+  ad=5.782e+11p pd=5.13e+06u as=0p ps=0u
M1010 a_410_58# a_811_379# a_231_132# VPB pshort w=840000u l=180000u
+  ad=4.83e+11p pd=2.83e+06u as=0p ps=0u
M1011 a_1852_374# B a_811_379# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.688e+11p ps=2.32e+06u
M1012 a_231_132# CI VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_811_379# a_879_55# a_1660_374# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2342_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1015 VPWR a_83_21# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1016 a_231_132# a_1023_379# a_410_58# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_83_21# a_811_379# a_644_104# VPB pshort w=840000u l=180000u
+  ad=7.392e+11p pd=3.44e+06u as=0p ps=0u
M1018 VGND A a_1852_374# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_879_55# a_1023_379# a_410_58# VPB pshort w=840000u l=180000u
+  ad=3.742e+11p pd=2.95e+06u as=0p ps=0u
M1020 a_644_104# a_1023_379# a_83_21# VNB nlowvt w=640000u l=150000u
+  ad=4.1745e+11p pd=3.87e+06u as=0p ps=0u
M1021 VPWR B a_879_55# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_2342_48# a_1660_374# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B a_879_55# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1660_374# B a_811_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_644_104# a_231_132# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_83_21# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1027 a_1852_374# B a_1023_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_231_132# a_1023_379# a_83_21# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2342_48# a_1660_374# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_1852_374# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2342_48# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fah_2 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_416_392# A VGND VNB nlowvt w=640000u l=150000u
+  ad=4.247e+11p pd=4.22e+06u as=1.82425e+12p ps=1.593e+07u
M1001 COUT a_1454_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=2.404e+12p ps=1.999e+07u
M1002 a_852_424# a_481_379# a_117_368# VPB pshort w=840000u l=180000u
+  ad=1.1046e+12p pd=4.31e+06u as=6.58e+11p ps=5.31e+06u
M1003 a_517_424# B a_416_392# VNB nlowvt w=640000u l=150000u
+  ad=3.904e+11p pd=2.5e+06u as=0p ps=0u
M1004 a_852_424# B a_117_368# VNB nlowvt w=640000u l=150000u
+  ad=4.448e+11p pd=2.67e+06u as=7.401e+11p ps=4.99e+06u
M1005 a_117_368# a_481_379# a_517_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_1454_424# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_1898_424# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 a_1898_424# a_852_424# a_1692_424# VNB nlowvt w=640000u l=150000u
+  ad=4.729e+11p pd=2.9e+06u as=6.112e+11p ps=4.47e+06u
M1009 SUM a_1898_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_1692_424# a_2055_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.12e+06u
M1011 COUT a_1454_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 VGND A a_81_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.272e+11p ps=1.99e+06u
M1013 a_1454_424# a_852_424# a_481_379# VNB nlowvt w=640000u l=150000u
+  ad=5.6e+11p pd=3.03e+06u as=2.33e+11p ps=2.13e+06u
M1014 a_416_392# B a_852_424# VPB pshort w=840000u l=180000u
+  ad=5.398e+11p pd=4.87e+06u as=0p ps=0u
M1015 a_1692_424# a_517_424# a_1454_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1898_424# a_517_424# a_1692_424# VPB pshort w=840000u l=180000u
+  ad=5.082e+11p pd=2.89e+06u as=9.84e+11p ps=5.92e+06u
M1017 a_1692_424# CI VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1898_424# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.146e+11p ps=2.06e+06u
M1019 a_416_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1692_424# a_2055_424# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.642e+11p ps=3.01e+06u
M1021 a_1454_424# a_517_424# a_481_379# VPB pshort w=840000u l=180000u
+  ad=8.484e+11p pd=3.7e+06u as=3.654e+11p ps=2.93e+06u
M1022 a_2055_424# a_852_424# a_1898_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1692_424# CI VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_117_368# a_81_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_481_379# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1692_424# a_852_424# a_1454_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_416_392# a_481_379# a_852_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_2055_424# a_517_424# a_1898_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A a_81_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1030 a_517_424# a_481_379# a_416_392# VPB pshort w=840000u l=180000u
+  ad=7.434e+11p pd=3.45e+06u as=0p ps=0u
M1031 SUM a_1898_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_117_368# B a_517_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_481_379# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_117_368# a_81_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_1454_424# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fah_4 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_1268_379# a_531_362# a_586_257# VPB pshort w=840000u l=180000u
+  ad=3.486e+11p pd=2.51e+06u as=3.7495e+11p ps=2.95e+06u
M1001 a_1183_102# a_536_114# a_1278_102# VPB pshort w=840000u l=180000u
+  ad=3.63125e+11p pd=2.94e+06u as=6.468e+11p ps=3.22e+06u
M1002 VGND a_1278_102# SUM VNB nlowvt w=740000u l=150000u
+  ad=3.15805e+12p pd=2.382e+07u as=4.144e+11p ps=4.08e+06u
M1003 a_430_362# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=5.782e+11p pd=5.13e+06u as=4.54925e+12p ps=2.931e+07u
M1004 a_1378_125# a_536_114# a_1268_379# VPB pshort w=840000u l=180000u
+  ad=7.049e+11p pd=5.6e+06u as=0p ps=0u
M1005 VPWR A a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1006 a_200_74# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.337e+11p pd=5.7e+06u as=0p ps=0u
M1007 a_430_362# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.026e+11p pd=3.94e+06u as=0p ps=0u
M1008 COUT a_1268_379# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1009 COUT a_1268_379# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1010 a_586_257# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_1268_379# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 SUM a_1278_102# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=0p ps=0u
M1013 VPWR a_1278_102# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_1268_379# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_1278_102# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_1378_125# a_1183_102# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND CI a_1378_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.616e+11p ps=3.69e+06u
M1018 a_536_114# B a_430_362# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1019 a_200_74# a_586_257# a_531_362# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1020 VGND a_1378_125# a_1183_102# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.4305e+11p ps=3.95e+06u
M1021 a_1278_102# a_531_362# a_1183_102# VNB nlowvt w=640000u l=150000u
+  ad=2.44125e+11p pd=2.21e+06u as=0p ps=0u
M1022 COUT a_1268_379# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_536_114# B a_200_74# VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1024 VPWR a_1268_379# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_586_257# B VGND VNB nlowvt w=740000u l=150000u
+  ad=5.59925e+11p pd=5.19e+06u as=0p ps=0u
M1026 a_586_257# a_536_114# a_1268_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.3685e+11p ps=2.18e+06u
M1027 a_531_362# B a_200_74# VNB nlowvt w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=4.268e+11p ps=4.01e+06u
M1028 SUM a_1278_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_430_362# a_586_257# a_536_114# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_200_74# a_586_257# a_536_114# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_1278_102# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 SUM a_1278_102# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_531_362# B a_430_362# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR CI a_1378_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_430_362# a_586_257# a_531_362# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 COUT a_1268_379# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND A a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1038 a_200_74# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_1268_379# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1378_125# a_536_114# a_1278_102# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1268_379# a_531_362# a_1378_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 SUM a_1278_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1278_102# a_531_362# a_1378_125# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 VGND a_1857_368# a_1967_384# VNB nlowvt w=640000u l=150000u
+  ad=1.989e+12p pd=1.212e+07u as=2.808e+11p ps=2.29e+06u
M1001 COUT a_430_418# a_1200_368# VNB nlowvt w=640000u l=150000u
+  ad=9.056e+11p pd=4.11e+06u as=1.792e+11p ps=1.84e+06u
M1002 a_1857_368# CIN VGND VNB nlowvt w=740000u l=150000u
+  ad=2.33e+11p pd=2.13e+06u as=0p ps=0u
M1003 a_1857_368# CIN VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=7.3255e+11p pd=5.84e+06u as=2.058e+12p ps=1.28e+07u
M1004 a_608_74# B a_28_74# VNB nlowvt w=640000u l=150000u
+  ad=3.40325e+11p pd=2.79e+06u as=3.901e+11p ps=3.89e+06u
M1005 a_1200_368# a_492_48# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.85e+11p pd=2.81e+06u as=0p ps=0u
M1006 a_259_368# a_492_48# a_430_418# VPB pshort w=840000u l=180000u
+  ad=5.404e+11p pd=4.86e+06u as=5.082e+11p ps=4.57e+06u
M1007 a_28_74# a_492_48# a_608_74# VPB pshort w=840000u l=180000u
+  ad=7.63e+11p pd=5.55e+06u as=3.32325e+11p ps=2.78e+06u
M1008 a_430_418# B a_28_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_259_368# a_28_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=5.088e+11p pd=4.15e+06u as=0p ps=0u
M1010 a_1967_384# a_430_418# a_2004_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.088e+11p ps=2.87e+06u
M1011 SUM a_2004_136# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1012 a_2004_136# a_608_74# a_1967_384# VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=5.152e+11p ps=4.8e+06u
M1013 a_1598_400# a_430_418# COUT VPB pshort w=840000u l=180000u
+  ad=3.98e+11p pd=2.82e+06u as=1.029e+12p ps=4.13e+06u
M1014 a_28_74# a_492_48# a_430_418# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.648e+11p ps=3.7e+06u
M1015 a_1857_368# a_430_418# a_2004_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_492_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.22e+11p ps=2.08e+06u
M1017 VGND A a_28_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_2004_136# a_608_74# a_1857_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 COUT a_608_74# a_1200_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND CIN a_1598_400# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1021 SUM a_2004_136# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_608_74# B a_259_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1598_400# a_608_74# COUT VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_259_368# a_28_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_259_368# a_492_48# a_608_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1200_368# a_492_48# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR CIN a_1598_400# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1857_368# a_1967_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_430_418# B a_259_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR B a_492_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
M1000 a_372_365# a_336_263# a_244_368# VPB pshort w=840000u l=180000u
+  ad=3.276e+11p pd=2.46e+06u as=6.6325e+11p ps=5.18e+06u
M1001 a_1026_389# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.43e+11p pd=2.71e+06u as=1.6192e+12p ps=1.192e+07u
M1002 a_244_368# a_27_100# VGND VNB nlowvt w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=1.579e+12p ps=1.063e+07u
M1003 a_374_120# a_336_263# a_244_368# VNB nlowvt w=640000u l=150000u
+  ad=3.0045e+11p pd=2.29e+06u as=0p ps=0u
M1004 a_1609_368# CI VGND VNB nlowvt w=740000u l=150000u
+  ad=2.589e+11p pd=2.2e+06u as=0p ps=0u
M1005 VPWR CI a_1264_421# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=9.136e+11p ps=4.08e+06u
M1006 a_1609_368# CI VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=5.488e+11p pd=5.04e+06u as=0p ps=0u
M1007 a_1744_94# a_372_365# a_1719_368# VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=6.707e+11p ps=5.55e+06u
M1008 a_27_100# B a_372_365# VPB pshort w=840000u l=180000u
+  ad=5.404e+11p pd=5.02e+06u as=0p ps=0u
M1009 SUM a_1744_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 a_1609_368# a_374_120# a_1744_94# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_374_120# a_336_263# a_27_100# VPB pshort w=840000u l=180000u
+  ad=3.976e+11p pd=2.8e+06u as=0p ps=0u
M1012 COUT_N a_374_120# a_1026_389# VPB pshort w=840000u l=180000u
+  ad=3.99e+11p pd=2.63e+06u as=0p ps=0u
M1013 a_27_100# B a_374_120# VNB nlowvt w=640000u l=150000u
+  ad=3.965e+11p pd=3.91e+06u as=0p ps=0u
M1014 VGND A a_27_100# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_244_368# B a_372_365# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.912e+11p ps=2.19e+06u
M1016 COUT_N a_372_365# a_1026_389# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=2.4e+06u as=4.992e+11p ps=2.84e+06u
M1017 VGND a_1609_368# a_1719_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.264e+11p ps=2.3e+06u
M1018 a_1264_421# a_374_120# COUT_N VNB nlowvt w=640000u l=150000u
+  ad=3.52e+11p pd=2.38e+06u as=0p ps=0u
M1019 a_244_368# B a_374_120# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_27_100# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_244_368# a_27_100# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1719_368# a_374_120# a_1744_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.224e+11p ps=2.6e+06u
M1023 a_1264_421# a_372_365# COUT_N VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B a_336_263# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=2.74e+06u
M1025 VGND CI a_1264_421# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1744_94# a_372_365# a_1609_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR B a_336_263# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1028 VPWR a_1609_368# a_1719_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 SUM a_1744_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1030 a_372_365# a_336_263# a_27_100# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1026_389# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fill_1 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fill_2 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fill_4 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fill_8 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fill_diode_2 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fill_diode_4 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fill_diode_8 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ha_1 A B VGND VNB VPB VPWR COUT SUM
M1000 VPWR A a_239_294# VPB pshort w=840000u l=180000u
+  ad=1.6456e+12p pd=9.84e+06u as=2.268e+11p ps=2.22e+06u
M1001 a_695_119# B a_239_294# VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.824e+11p ps=1.85e+06u
M1002 VPWR A a_389_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.9e+11p ps=2.78e+06u
M1003 a_389_392# B a_83_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.13e+11p ps=2.65e+06u
M1004 COUT a_239_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=6.95225e+11p ps=6.36e+06u
M1005 VPWR a_83_260# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1006 a_83_260# a_239_294# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_305_130# a_239_294# a_83_260# VNB nlowvt w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=1.726e+11p ps=1.85e+06u
M1008 COUT a_239_294# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1009 VGND B a_305_130# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_695_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_83_260# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1012 a_239_294# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_305_130# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ha_2 A B VGND VNB VPB VPWR COUT SUM
M1000 COUT a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.01665e+12p ps=1.023e+07u
M1001 a_278_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.083e+11p pd=4.09e+06u as=0p ps=0u
M1002 SUM a_394_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.9664e+12p ps=1.448e+07u
M1003 VPWR a_394_388# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 SUM a_394_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=0p ps=0u
M1005 a_310_388# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1006 COUT a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1007 VGND B a_278_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_74# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1010 a_394_388# B a_310_388# VPB pshort w=1e+06u l=180000u
+  ad=9.6e+11p pd=3.92e+06u as=0p ps=0u
M1011 VPWR a_27_74# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_394_388# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_27_74# a_394_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1015 VPWR A a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_114_74# B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_278_74# a_27_74# a_394_388# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.01625e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ha_4 A B VGND VNB VPB VPWR COUT SUM
M1000 a_435_99# B a_707_119# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=5.856e+11p ps=5.67e+06u
M1001 a_297_392# a_435_99# VPWR VPB pshort w=840000u l=180000u
+  ad=4.968e+11p pd=4.76e+06u as=2.6878e+12p ps=2.354e+07u
M1002 VGND B a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=1.6734e+12p pd=1.601e+07u as=7.744e+11p ps=7.54e+06u
M1003 a_707_119# B a_435_99# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_707_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_297_392# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.069e+11p ps=4.33e+06u
M1006 VPWR a_435_99# a_297_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_125# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_435_99# B VPWR VPB pshort w=840000u l=180000u
+  ad=7.46425e+11p pd=5.89e+06u as=0p ps=0u
M1009 COUT a_435_99# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=7.84e+11p pd=5.88e+06u as=0p ps=0u
M1010 VGND a_435_99# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1011 a_707_119# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_435_99# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_125# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_435_99# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 SUM a_297_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=8.1e+11p ps=7.62e+06u
M1017 a_27_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 COUT a_435_99# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_297_392# B a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_435_99# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_392# B a_297_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_297_392# a_435_99# a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=0p ps=0u
M1024 SUM a_297_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=8.96e+11p pd=6.08e+06u as=0p ps=0u
M1025 VPWR B a_435_99# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 SUM a_297_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_297_392# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_125# a_435_99# a_297_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_435_99# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_297_392# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 SUM a_297_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 COUT a_435_99# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 COUT a_435_99# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR A a_435_99# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_297_392# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__inv_1 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.627e+11p ps=2.19e+06u
M1001 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=3.696e+11p ps=2.9e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__inv_16 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=1.6576e+12p pd=1.632e+07u as=2.2718e+12p ps=1.946e+07u
M1001 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.4528e+12p pd=2.23e+07u as=3.1584e+12p ps=2.58e+07u
M1005 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__inv_2 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=6.048e+11p ps=5.56e+06u
M1001 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=4.218e+11p ps=4.1e+06u
M1003 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__inv_4 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.296e+11p ps=8.38e+06u
M1001 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=6.882e+11p pd=6.3e+06u as=4.44e+11p ps=4.16e+06u
M1003 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__inv_8 A VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=1.2025e+12p pd=1.065e+07u as=8.288e+11p ps=8.16e+06u
M1001 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=1.7024e+12p ps=1.424e+07u
M1003 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__maj3_1 A B C VGND VNB VPB VPWR X
M1000 a_601_384# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=7.15e+11p ps=5.61e+06u
M1001 VPWR a_84_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1002 VGND a_84_74# X VNB nlowvt w=740000u l=150000u
+  ad=5.466e+11p pd=4.39e+06u as=2.081e+11p ps=2.05e+06u
M1003 a_84_74# C a_601_384# VPB pshort w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 a_84_74# B a_223_120# VNB nlowvt w=640000u l=150000u
+  ad=4.177e+11p pd=4.01e+06u as=1.536e+11p ps=1.76e+06u
M1005 a_595_136# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1006 a_229_384# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 VGND C a_403_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1008 a_84_74# C a_595_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_409_384# B a_84_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1010 a_84_74# B a_229_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_223_120# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C a_409_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_403_136# B a_84_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__maj3_2 A B C VGND VNB VPB VPWR X
M1000 a_396_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.43375e+11p pd=2.86e+06u as=1.495e+12p ps=9.5e+06u
M1001 VPWR C a_587_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1002 a_577_74# B a_87_264# VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=4.181e+11p ps=4.09e+06u
M1003 VGND C a_577_74# VNB nlowvt w=740000u l=150000u
+  ad=1.2062e+12p pd=7.7e+06u as=0p ps=0u
M1004 VPWR a_87_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1005 X a_87_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_793_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 a_87_264# B a_396_368# VPB pshort w=1e+06u l=180000u
+  ad=5.5e+11p pd=5.1e+06u as=0p ps=0u
M1008 a_413_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1009 a_87_264# B a_413_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_587_347# B a_87_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_87_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1012 a_793_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1013 a_87_264# C a_793_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_87_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_87_264# C a_793_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__maj3_4 A B C VGND VNB VPB VPWR X
M1000 a_222_392# B a_504_125# VNB nlowvt w=640000u l=150000u
+  ad=5.376e+11p pd=5.52e+06u as=5.41775e+11p ps=4.6e+06u
M1001 X a_222_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=1.2479e+12p ps=1.196e+07u
M1002 a_908_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=1.971e+12p ps=1.647e+07u
M1003 a_222_392# C a_906_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.45475e+11p ps=4.25e+06u
M1004 a_222_392# B a_122_392# VPB pshort w=1e+06u l=180000u
+  ad=8.6e+11p pd=7.72e+06u as=5.9e+11p ps=5.18e+06u
M1005 a_222_392# C a_908_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_906_78# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_122_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_122_392# B a_222_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_122_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_504_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_906_78# C a_222_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A a_906_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_908_392# C a_222_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A a_908_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_114_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.7375e+11p ps=4.61e+06u
M1016 X a_222_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1017 a_114_125# B a_222_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_504_125# C VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_222_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_222_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_114_125# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_222_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_222_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_222_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_222_392# B a_114_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_504_125# B a_222_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_222_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_504_392# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1029 VPWR C a_504_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_504_392# B a_222_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_222_392# B a_504_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2_1 A0 A1 S VGND VNB VPB VPWR X
M1000 a_304_74# A0 a_226_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=7.85e+11p ps=3.57e+06u
M1001 X a_304_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=8.226e+11p ps=5.83e+06u
M1002 a_443_74# A0 a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=3.1e+06u as=4.033e+11p ps=2.57e+06u
M1003 VPWR S a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1004 VPWR a_27_112# a_527_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.9e+11p ps=2.78e+06u
M1005 a_527_368# A1 a_304_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND S a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=7.0725e+11p pd=4.91e+06u as=1.5675e+11p ps=1.67e+06u
M1007 a_304_74# A1 a_226_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1008 a_226_74# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_112# a_443_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_304_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1011 a_226_368# S VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2_2 A0 A1 S VGND VNB VPB VPWR X
M1000 a_119_368# A0 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=5.6e+11p ps=5.12e+06u
M1001 a_209_368# A1 a_119_368# VPB pshort w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1002 a_119_368# A0 a_38_74# VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=2.63e+06u as=4.292e+11p ps=4.12e+06u
M1003 X a_119_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=9.4915e+11p ps=7.09e+06u
M1004 a_38_74# a_459_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_209_368# a_459_48# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.133e+12p ps=8.62e+06u
M1006 a_270_74# A1 a_119_368# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1007 VPWR S a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR S a_459_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 VGND S a_270_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_119_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1011 VPWR a_119_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND S a_459_48# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 VGND a_119_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2_4 A0 A1 S VGND VNB VPB VPWR X
M1000 X a_193_241# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.06535e+12p pd=6.79e+06u as=2.35648e+12p ps=1.609e+07u
M1001 a_709_119# S VGND VNB nlowvt w=640000u l=150000u
+  ad=4.224e+11p pd=3.88e+06u as=1.76805e+12p ps=1.249e+07u
M1002 VGND S a_27_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1003 a_937_119# a_27_368# VGND VNB nlowvt w=640000u l=150000u
+  ad=3.712e+11p pd=3.72e+06u as=0p ps=0u
M1004 X a_193_241# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_939_391# A1 a_193_241# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=9.25e+11p ps=7.85e+06u
M1006 X a_193_241# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=0p ps=0u
M1007 VGND a_27_368# a_937_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_193_241# A1 a_939_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR S a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1010 a_725_391# S VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1011 a_725_391# A0 a_193_241# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_193_241# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR S a_725_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_193_241# A1 a_709_119# VNB nlowvt w=640000u l=150000u
+  ad=9.216e+11p pd=6.72e+06u as=0p ps=0u
M1015 a_939_391# a_27_368# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_193_241# A0 a_725_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_937_119# A0 a_193_241# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_27_368# a_939_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_193_241# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_193_241# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_193_241# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_193_241# A0 a_937_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_193_241# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND S a_709_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_709_119# A1 a_193_241# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
M1000 Y A0 a_426_74# VNB nlowvt w=740000u l=150000u
+  ad=5.217e+11p pd=2.89e+06u as=1.776e+11p ps=1.96e+06u
M1001 a_426_74# a_114_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.6755e+11p ps=3.99e+06u
M1002 VPWR S a_223_368# VPB pshort w=1.12e+06u l=180000u
+  ad=5.292e+11p pd=5e+06u as=5.936e+11p ps=5.54e+06u
M1003 a_402_368# a_114_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=0p ps=0u
M1004 a_225_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=0p ps=0u
M1005 Y A0 a_223_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 a_402_368# A1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_114_74# S VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1008 VGND S a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_114_74# S VPWR VPB pshort w=840000u l=180000u
+  ad=2.184e+11p pd=2.2e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
M1000 VPWR a_922_72# a_343_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.58023e+12p pd=1.017e+07u as=1.0304e+12p ps=6.32e+06u
M1001 VGND a_922_72# a_115_74# VNB nlowvt w=740000u l=150000u
+  ad=1.10195e+12p pd=8.18e+06u as=5.18e+11p ps=4.36e+06u
M1002 Y A0 a_121_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1312e+12p pd=8.74e+06u as=6.496e+11p ps=5.64e+06u
M1003 Y A1 a_343_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_922_72# S VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1005 a_337_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=7.8555e+11p pd=5.15e+06u as=8.4255e+11p ps=6.93e+06u
M1006 a_121_368# S VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR S a_121_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_115_74# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_922_72# S VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1010 a_337_74# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_121_368# A0 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_343_368# a_922_72# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND S a_337_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_343_368# A1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_337_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A0 a_115_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_115_74# a_922_72# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
M1000 Y A1 a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=1.0767e+12p pd=1.031e+07u as=8.917e+11p ps=8.33e+06u
M1001 a_481_368# A0 Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.3104e+12p pd=1.13e+07u as=1.6576e+12p ps=1.416e+07u
M1002 VPWR a_1030_268# a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.387e+12p pd=1.732e+07u as=1.2992e+12p ps=1.128e+07u
M1003 a_481_368# S VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR S a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_114_85# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR S a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_475_85# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=8.806e+11p pd=8.3e+06u as=0p ps=0u
M1008 a_119_368# A1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_114_85# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.795e+12p ps=1.331e+07u
M1011 a_119_368# A1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_119_368# a_1030_268# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_475_85# a_1030_268# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_1030_268# a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A0 a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_114_85# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A0 a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_481_368# A0 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1030_268# a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_119_368# a_1030_268# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_114_85# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A1 a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1030_268# S VGND VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1025 VGND S a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_1030_268# a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1030_268# S VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1028 VGND S a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_475_85# a_1030_268# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A0 a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A0 a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_481_368# S VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR S a_1030_268# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_475_85# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_540_341# VPB pshort w=1e+06u l=180000u
+  ad=1.87058e+12p pd=1.254e+07u as=3.3e+11p ps=2.66e+06u
M1001 VGND A1 a_450_74# VNB nlowvt w=640000u l=150000u
+  ad=1.2058e+12p pd=9.01e+06u as=4.8e+11p ps=2.78e+06u
M1002 a_766_341# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.6525e+11p pd=3.11e+06u as=0p ps=0u
M1003 a_979_74# S0 a_846_74# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=7.84075e+11p ps=5.5e+06u
M1004 a_1338_125# S1 a_846_74# VNB nlowvt w=640000u l=150000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1005 a_1068_387# a_27_74# a_846_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=1.155e+12p ps=6.31e+06u
M1006 a_846_74# a_1396_99# a_1338_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1007 a_1338_125# S1 a_342_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.5e+11p ps=5.1e+06u
M1008 a_846_74# S0 a_766_341# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR S0 a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1010 a_342_74# S0 a_258_341# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.8e+11p ps=3.56e+06u
M1011 VGND S1 a_1396_99# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1012 VPWR A3 a_1068_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_540_341# a_27_74# a_342_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_264_74# A0 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1015 a_342_74# a_27_74# a_264_74# VNB nlowvt w=640000u l=150000u
+  ad=4.32e+11p pd=3.91e+06u as=0p ps=0u
M1016 VPWR S1 a_1396_99# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1017 X a_1338_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1018 X a_1338_125# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1019 a_450_74# S0 a_342_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_258_341# A0 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND S0 a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1022 a_846_74# a_27_74# a_768_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1023 a_768_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_342_74# a_1396_99# a_1338_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A3 a_979_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 VGND S0 a_31_94# VNB nlowvt w=640000u l=150000u
+  ad=1.6907e+12p pd=1.216e+07u as=1.824e+11p ps=1.85e+06u
M1001 VPWR S0 a_31_94# VPB pshort w=1e+06u l=180000u
+  ad=2.256e+12p pd=1.486e+07u as=2.8e+11p ps=2.56e+06u
M1002 a_1155_392# S0 a_909_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=7.85e+11p ps=5.57e+06u
M1003 a_1429_74# S1 a_333_74# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=8.45e+11p ps=5.69e+06u
M1004 a_1047_74# a_31_94# a_909_74# VNB nlowvt w=740000u l=150000u
+  ad=5.772e+11p pd=3.04e+06u as=6.068e+11p ps=4.6e+06u
M1005 a_909_74# a_31_94# a_843_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.9e+11p ps=3.38e+06u
M1006 a_909_74# a_1500_94# a_1429_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_333_74# a_1500_94# a_1429_74# VNB nlowvt w=740000u l=150000u
+  ad=7.437e+11p pd=4.97e+06u as=3.0295e+11p ps=2.65e+06u
M1008 a_621_392# S0 a_333_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1009 VGND S1 a_1500_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.76725e+11p ps=2.15e+06u
M1010 a_1429_74# S1 a_909_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_333_74# S0 a_255_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1012 VGND A2 a_1047_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_255_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_507_74# a_31_94# a_333_74# VNB nlowvt w=740000u l=150000u
+  ad=5.772e+11p pd=3.04e+06u as=0p ps=0u
M1015 X a_1429_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1016 a_909_74# S0 a_831_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1017 VPWR A0 a_621_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_843_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A2 a_1155_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_831_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_1429_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_1429_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1023 a_333_74# a_31_94# a_267_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=8.7e+11p ps=3.74e+06u
M1024 VGND A0 a_507_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_1429_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_267_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR S1 a_1500_94# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.1e+11p ps=2.82e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 a_509_392# S0 a_299_392# VPB pshort w=1e+06u l=180000u
+  ad=1.19e+12p pd=1.038e+07u as=6.15e+11p ps=5.23e+06u
M1001 a_1468_377# S0 a_1191_121# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=1.15e+12p ps=1.03e+07u
M1002 a_1278_121# a_758_306# a_1191_121# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=9.2755e+11p ps=8.21e+06u
M1003 a_119_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=3.48045e+12p ps=2.828e+07u
M1004 VPWR A1 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1288_377# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1006 a_1191_121# a_758_306# a_1278_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A0 a_299_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1191_121# S0 a_1468_377# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_509_392# S0 a_114_126# VNB nlowvt w=640000u l=150000u
+  ad=8.5705e+11p pd=8.11e+06u as=3.872e+11p ps=3.77e+06u
M1010 X a_2199_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1011 a_299_392# A0 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1450_121# S0 a_1191_121# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1013 VPWR S0 a_758_306# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1014 VGND S1 a_2489_347# VNB nlowvt w=740000u l=150000u
+  ad=2.4642e+12p pd=2.151e+07u as=2.109e+11p ps=2.05e+06u
M1015 a_2199_74# a_2489_347# a_509_392# VNB nlowvt w=640000u l=150000u
+  ad=8.576e+11p pd=6.52e+06u as=0p ps=0u
M1016 VGND S0 a_758_306# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_1191_121# S1 a_2199_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1450_121# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_2199_74# S1 a_1191_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_2199_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1021 a_1278_121# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_299_126# A0 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1023 VGND A0 a_299_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A3 a_1288_377# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A1 a_114_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_2199_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_2199_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1191_121# a_2489_347# a_2199_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=9.3e+11p ps=7.86e+06u
M1029 a_2199_74# a_2489_347# a_1191_121# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_2199_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A3 a_1450_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2199_74# S1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_114_126# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_2199_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_2199_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1468_377# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_509_392# S1 a_2199_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR A2 a_1468_377# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_299_126# a_758_306# a_509_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND A2 a_1278_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1191_121# S0 a_1450_121# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_299_392# S0 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_509_392# a_758_306# a_299_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR S1 a_2489_347# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.528e+11p ps=2.87e+06u
M1045 a_119_392# a_758_306# a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1288_377# a_758_306# a_1191_121# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_114_126# S0 a_509_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_509_392# a_2489_347# a_2199_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_509_392# a_758_306# a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_1191_121# a_758_306# a_1288_377# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1051 X a_2199_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand2_1 A B VGND VNB VPB VPWR Y
M1000 Y A a_117_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.776e+11p ps=1.96e+06u
M1001 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=6.048e+11p ps=5.56e+06u
M1002 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand2_2 A B VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.408e+11p ps=8.4e+06u
M1001 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=6.438e+11p ps=6.18e+06u
M1003 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.442e+11p ps=2.14e+06u
M1006 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand2_4 A B VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.0472e+12p pd=8.59e+06u as=2.6824e+12p ps=9.27e+06u
M1001 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=5.365e+11p pd=4.41e+06u as=1.1581e+12p ps=1.053e+07u
M1003 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1005 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand2_8 A B VGND VNB VPB VPWR Y
M1000 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=1.0656e+12p pd=8.8e+06u as=2.14795e+12p ps=1.918e+07u
M1001 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.288e+11p ps=8.16e+06u
M1004 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=5.0008e+12p pd=2.237e+07u as=1.3216e+12p ps=1.132e+07u
M1007 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand2b_1 A_N B VGND VNB VPB VPWR Y
M1000 Y a_27_112# a_269_74# VNB nlowvt w=740000u l=150000u
+  ad=3.182e+11p pd=2.34e+06u as=1.776e+11p ps=1.96e+06u
M1001 a_269_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.4825e+11p ps=2.73e+06u
M1002 VPWR A_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=8.47e+11p pd=6.03e+06u as=2.352e+11p ps=2.24e+06u
M1003 VGND A_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1004 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.584e+11p pd=2.88e+06u as=0p ps=0u
M1005 VPWR a_27_112# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand2b_2 A_N B VGND VNB VPB VPWR Y
M1000 Y a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.5068e+12p ps=9.46e+06u
M1001 VPWR a_27_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND B a_242_74# VNB nlowvt w=740000u l=150000u
+  ad=3.7765e+11p pd=3.86e+06u as=6.2445e+11p ps=6.14e+06u
M1003 VPWR A_N a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1004 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_27_74# a_242_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1007 a_242_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A_N a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1009 a_242_74# a_27_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand2b_4 A_N B VGND VNB VPB VPWR Y
M1000 Y a_31_74# a_243_74# VNB nlowvt w=740000u l=150000u
+  ad=5.143e+11p pd=4.35e+06u as=1.0434e+12p ps=1.022e+07u
M1001 a_243_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.0286e+12p ps=7.22e+06u
M1002 a_31_74# A_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=2.9792e+12p ps=1.407e+07u
M1003 VGND B a_243_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.0528e+12p pd=6.36e+06u as=0p ps=0u
M1005 VPWR A_N a_31_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_31_74# a_243_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_243_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_243_74# a_31_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B a_243_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A_N a_31_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 VPWR a_31_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_243_74# a_31_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_31_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand3_1 A B C VGND VNB VPB VPWR Y
M1000 Y A a_233_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=3.108e+11p ps=2.32e+06u
M1001 a_233_74# B a_155_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1002 a_155_74# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1003 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=8.4e+11p ps=5.98e+06u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand3_2 A B C VGND VNB VPB VPWR Y
M1000 a_27_74# C VGND VNB nlowvt w=740000u l=150000u
+  ad=6.068e+11p pd=6.08e+06u as=2.072e+11p ps=2.04e+06u
M1001 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.3384e+12p pd=1.135e+07u as=9.128e+11p ps=8.35e+06u
M1002 a_283_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=7.123e+11p pd=5.5e+06u as=2.072e+11p ps=2.04e+06u
M1003 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_283_74# B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# B a_283_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A a_283_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand3_4 A B C VGND VNB VPB VPWR Y
M1000 a_456_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=8.288e+11p pd=8.16e+06u as=6.142e+11p ps=6.1e+06u
M1001 VGND C a_456_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_82# B a_456_82# VNB nlowvt w=740000u l=150000u
+  ad=1.0121e+12p pd=1.018e+07u as=0p ps=0u
M1003 a_456_82# B a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.4896e+12p pd=9.38e+06u as=3.5896e+12p ps=1.537e+07u
M1005 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1008 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_456_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_82# B a_456_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_456_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_82# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_456_82# B a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_82# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand3b_1 A_N B C VGND VNB VPB VPWR Y
M1000 Y a_27_116# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=8.47e+11p ps=6.03e+06u
M1001 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y a_27_116# a_347_78# VNB nlowvt w=740000u l=150000u
+  ad=3.404e+11p pd=2.4e+06u as=2.886e+11p ps=2.26e+06u
M1003 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A_N a_27_116# VNB nlowvt w=550000u l=150000u
+  ad=4.4825e+11p pd=2.73e+06u as=1.5675e+11p ps=1.67e+06u
M1005 VPWR A_N a_27_116# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 a_269_78# C VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1007 a_347_78# B a_269_78# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand3b_2 A_N B C VGND VNB VPB VPWR Y
M1000 VPWR A_N a_27_94# VPB pshort w=1e+06u l=180000u
+  ad=1.5646e+12p pd=1.177e+07u as=2.8e+11p ps=2.56e+06u
M1001 a_206_74# C VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=4.2745e+11p ps=4.18e+06u
M1002 VGND A_N a_27_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1003 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.0248e+12p ps=8.55e+06u
M1004 Y a_27_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_27_94# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_27_94# a_403_54# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.1145e+11p ps=7.38e+06u
M1007 a_403_54# a_27_94# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C a_206_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_206_74# B a_403_54# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_403_54# B a_206_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand3b_4 A_N B C VGND VNB VPB VPWR Y
M1000 VGND A_N a_89_172# VNB nlowvt w=740000u l=150000u
+  ad=1.1492e+12p pd=8.02e+06u as=1.9515e+11p ps=2.05e+06u
M1001 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=4.8426e+12p pd=1.966e+07u as=1.3328e+12p ps=9.1e+06u
M1002 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_744_74# B a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=1.0672e+12p pd=1.036e+07u as=8.806e+11p ps=8.3e+06u
M1004 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_744_74# a_89_172# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=4.13e+06u
M1006 a_297_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_744_74# B a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_89_172# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_89_172# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_297_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_89_172# a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_89_172# a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_297_82# B a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_297_82# B a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_89_172# A_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1018 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_744_74# a_89_172# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A_N a_89_172# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4_1 A B C D VGND VNB VPB VPWR Y
M1000 a_181_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.923e+11p ps=2.72e+06u
M1001 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.608e+11p pd=5.66e+06u as=1.1648e+12p ps=8.8e+06u
M1002 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_259_74# C a_181_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1004 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_373_74# B a_259_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1007 Y A a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=2.085e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4_2 A B C D VGND VNB VPB VPWR Y
M1000 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=2.1336e+12p pd=1.501e+07u as=1.2768e+12p ps=1.124e+07u
M1001 a_515_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=6.2875e+11p pd=6.24e+06u as=2.22e+11p ps=2.08e+06u
M1002 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=6.5035e+11p pd=6.28e+06u as=2.738e+11p ps=2.22e+06u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_515_74# B a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1008 a_304_74# C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A a_515_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND D a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# C a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_304_74# B a_515_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4_4 A B C D VGND VNB VPB VPWR Y
M1000 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=5.1016e+12p pd=2.031e+07u as=2.6544e+12p ps=1.37e+07u
M1001 a_554_74# C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=8.288e+11p pd=8.16e+06u as=1.13125e+12p ps=1.05e+07u
M1002 Y A a_923_74# VNB nlowvt w=740000u l=150000u
+  ad=5.328e+11p pd=4.4e+06u as=1.0147e+12p ps=1.022e+07u
M1003 a_923_74# B a_554_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_923_74# B a_554_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND D a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=6.66e+11p pd=4.76e+06u as=0p ps=0u
M1007 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# C a_554_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_554_74# C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_923_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A a_923_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_554_74# B a_923_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND D a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_74# C a_554_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_554_74# B a_923_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_923_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.239e+12p ps=8.97e+06u
M1001 VPWR a_27_112# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_443_74# B a_341_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=2.664e+11p ps=2.2e+06u
M1003 Y a_27_112# a_443_74# VNB nlowvt w=740000u l=150000u
+  ad=3.404e+11p pd=2.4e+06u as=0p ps=0u
M1004 VPWR A_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1005 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=2.696e+11p pd=2.26e+06u as=2.695e+11p ps=2.08e+06u
M1007 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_263_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1009 a_341_74# C a_263_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
M1000 a_719_123# C a_490_74# VNB nlowvt w=740000u l=150000u
+  ad=6.22175e+11p pd=6.14e+06u as=5.618e+11p ps=4.6e+06u
M1001 a_225_74# B a_490_74# VNB nlowvt w=740000u l=150000u
+  ad=6.01175e+11p pd=6.14e+06u as=0p ps=0u
M1002 a_225_74# a_27_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1003 a_719_123# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.946e+11p ps=3.93e+06u
M1004 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=2.3654e+12p ps=1.544e+07u
M1005 VGND D a_719_123# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_490_74# C a_719_123# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_490_74# B a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A_N a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1009 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A_N a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1011 Y a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_27_74# a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
M1000 a_656_74# C a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=8.399e+11p pd=8.19e+06u as=1.0287e+12p ps=1.022e+07u
M1001 VGND D a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=6.9465e+11p pd=6.36e+06u as=0p ps=0u
M1002 Y a_27_158# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.1168e+12p pd=1.274e+07u as=4.9266e+12p ps=2.188e+07u
M1003 a_225_74# B a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=1.01295e+12p pd=1.022e+07u as=0p ps=0u
M1004 VPWR a_27_158# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_225_74# a_27_158# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1006 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_1025_158# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1025_158# C a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_656_74# B a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_225_74# a_27_158# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1025_158# C a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1025_158# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND D a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_158# A_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1019 a_225_74# B a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_656_74# B a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A_N a_27_158# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A_N a_27_158# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.962e+11p ps=2.05e+06u
M1024 Y a_27_158# a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y a_27_158# a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_656_74# C a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
M1000 a_229_398# B_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5055e+11p pd=1.69e+06u as=5.10375e+11p ps=4.39e+06u
M1001 a_513_74# a_229_398# a_435_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=1.776e+11p ps=1.96e+06u
M1002 VGND A_N a_27_398# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.50975e+11p ps=1.67e+06u
M1003 VGND D a_627_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.108e+11p ps=2.32e+06u
M1004 VPWR a_27_398# Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.1844e+12p pd=8.46e+06u as=9.856e+11p ps=8.48e+06u
M1005 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_229_398# B_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1007 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_229_398# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_435_74# a_27_398# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.9585e+11p ps=2.05e+06u
M1010 VPWR A_N a_27_398# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1011 a_627_74# C a_513_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
M1000 Y a_231_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2544e+12p pd=1.12e+07u as=2.8737e+12p ps=1.85e+07u
M1001 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_373_74# a_231_74# a_678_74# VNB nlowvt w=740000u l=150000u
+  ad=8.504e+11p pd=6.86e+06u as=4.662e+11p ps=4.22e+06u
M1003 Y a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_231_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_231_74# B_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=5.278e+11p ps=4.3e+06u
M1006 a_886_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=0p ps=0u
M1007 VPWR a_27_368# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D a_886_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A_N a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1011 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_373_74# a_27_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.257e+11p ps=2.09e+06u
M1013 a_886_74# C a_678_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_678_74# a_231_74# a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_27_368# a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_231_74# B_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.8e+11p pd=2.76e+06u as=0p ps=0u
M1018 VGND A_N a_27_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1019 a_678_74# C a_886_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
M1000 VPWR a_27_114# Y VPB pshort w=1.12e+06u l=180000u
+  ad=3.64e+12p pd=3.044e+07u as=2.4752e+12p ps=2.234e+07u
M1001 a_374_74# a_27_114# Y VNB nlowvt w=740000u l=150000u
+  ad=1.0508e+12p pd=1.024e+07u as=4.921e+11p ps=4.29e+06u
M1002 Y a_27_114# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y a_27_114# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_828_74# a_232_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=9.53e+11p pd=8.52e+06u as=0p ps=0u
M1005 a_1229_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0434e+12p pd=1.022e+07u as=9.049e+11p ps=7.36e+06u
M1006 VPWR a_27_114# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_374_74# a_27_114# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_374_74# a_232_114# a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_232_114# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y a_27_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_232_114# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_828_74# a_232_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_114# A_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1016 VPWR A_N a_27_114# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_232_114# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A_N a_27_114# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1019 a_232_114# B_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1020 VPWR a_232_114# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_232_114# B_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=0p ps=0u
M1023 a_828_74# C a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR B_N a_232_114# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_828_74# C a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_374_74# a_232_114# a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y a_27_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1229_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1229_74# C a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1229_74# C a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2_1 A B VGND VNB VPB VPWR Y
M1000 a_119_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=3.136e+11p ps=2.8e+06u
M1001 Y B a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=2.072e+11p ps=2.04e+06u
M1003 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2_2 A B VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=5.254e+11p pd=4.38e+06u as=2.072e+11p ps=2.04e+06u
M1001 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B a_35_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=9.296e+11p ps=8.38e+06u
M1003 a_35_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A a_35_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 a_35_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2_4 A B VGND VNB VPB VPWR Y
M1000 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.6576e+12p ps=1.416e+07u
M1001 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=1.4874e+12p pd=8.46e+06u as=1.0656e+12p ps=5.84e+06u
M1003 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.608e+11p pd=5.66e+06u as=0p ps=0u
M1008 a_27_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2_8 A B VGND VNB VPB VPWR Y
M1000 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=2.1756e+12p pd=1.328e+07u as=1.4393e+12p ps=9.81e+06u
M1001 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+12p pd=2.536e+07u as=1.4336e+12p ps=1.152e+07u
M1002 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2656e+12p pd=1.122e+07u as=0p ps=0u
M1013 a_27_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2b_1 A B_N VGND VNB VPB VPWR Y
M1000 a_281_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=4.396e+11p ps=3.1e+06u
M1001 Y a_27_112# a_281_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=0p ps=0u
M1002 VGND a_27_112# Y VNB nlowvt w=740000u l=150000u
+  ad=5.6985e+11p pd=4.59e+06u as=2.627e+11p ps=2.19e+06u
M1003 VPWR B_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1004 VGND B_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.805e+11p ps=2.12e+06u
M1005 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2b_2 A B_N VGND VNB VPB VPWR Y
M1000 a_228_368# a_27_392# Y VPB pshort w=1.12e+06u l=180000u
+  ad=9.24e+11p pd=8.37e+06u as=3.024e+11p ps=2.78e+06u
M1001 VPWR A a_228_368# VPB pshort w=1.12e+06u l=180000u
+  ad=5.824e+11p pd=5.34e+06u as=0p ps=0u
M1002 a_228_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.884e+11p pd=4.28e+06u as=7.744e+11p ps=6.56e+06u
M1004 VPWR B_N a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1005 VGND B_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1006 VGND a_27_392# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_392# a_228_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2b_4 A B_N VGND VNB VPB VPWR Y
M1000 a_353_323# B_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=1.2838e+12p ps=1.087e+07u
M1001 a_353_323# B_N VGND VNB nlowvt w=740000u l=150000u
+  ad=5.18e+11p pd=2.88e+06u as=1.3489e+12p ps=8.29e+06u
M1002 VPWR B_N a_353_323# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1004 a_119_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2656e+12p pd=1.122e+07u as=0p ps=0u
M1005 VPWR A a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_353_323# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_119_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_353_323# a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1010 a_119_368# a_353_323# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y a_353_323# a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_368# a_353_323# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_353_323# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3_1 A B C VGND VNB VPB VPWR Y
M1000 Y C a_201_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=3.696e+11p ps=2.9e+06u
M1001 a_117_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=3.024e+11p ps=2.78e+06u
M1002 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=4.699e+11p ps=4.23e+06u
M1003 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_201_368# B a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3_2 A B C VGND VNB VPB VPWR Y
M1000 a_27_368# C Y VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=8.38e+06u as=3.584e+11p ps=2.88e+06u
M1001 a_309_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.384e+11p pd=5.62e+06u as=0p ps=0u
M1002 Y C a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_309_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.248e+11p ps=2.82e+06u
M1004 a_27_368# B a_309_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_309_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=9.176e+11p pd=5.44e+06u as=4.699e+11p ps=4.23e+06u
M1007 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3_4 A B C VGND VNB VPB VPWR Y
M1000 Y C a_298_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.786e+11p pd=6.44e+06u as=1.8418e+12p ps=1.279e+07u
M1001 Y C a_298_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=1.22935e+12p ps=9.25e+06u
M1003 a_27_368# B a_298_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.5176e+12p pd=1.391e+07u as=0p ps=0u
M1004 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_298_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.048e+11p ps=5.56e+06u
M1009 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_368# B a_298_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_298_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_298_368# C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_298_368# C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3b_1 A B C_N VGND VNB VPB VPWR Y
M1000 Y a_27_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.477e+11p pd=4.17e+06u as=5.8515e+11p ps=4.58e+06u
M1001 Y a_27_112# a_347_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=4.368e+11p ps=3.02e+06u
M1002 a_347_368# B a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.688e+11p ps=2.72e+06u
M1003 a_263_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.06e+11p ps=3.02e+06u
M1004 VGND C_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.695e+11p ps=2.08e+06u
M1005 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1007 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3b_2 A B C_N VGND VNB VPB VPWR Y
M1000 VGND a_27_392# Y VNB nlowvt w=740000u l=150000u
+  ad=1.6739e+12p pd=1.049e+07u as=6.697e+11p ps=6.25e+06u
M1001 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR C_N a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=8.91e+11p pd=8.13e+06u as=2.75e+11p ps=2.55e+06u
M1004 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_27_392# a_227_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=9.184e+11p ps=8.36e+06u
M1006 a_227_368# a_27_392# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_498_368# B a_227_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1008 VGND C_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1009 a_498_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_227_368# B a_498_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A a_498_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3b_4 A B C_N VGND VNB VPB VPWR Y
M1000 VGND a_468_264# Y VNB nlowvt w=740000u l=150000u
+  ad=2.0498e+12p pd=1.59e+07u as=1.3135e+12p ps=1.243e+07u
M1001 a_27_368# B a_129_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.5904e+12p pd=1.404e+07u as=1.2936e+12p ps=1.127e+07u
M1002 Y a_468_264# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1003 a_129_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.2838e+12p ps=1.087e+07u
M1004 Y a_468_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_368# a_468_264# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_129_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_368# B a_129_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_468_264# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_129_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_368# a_468_264# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_129_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_468_264# C_N VGND VNB nlowvt w=740000u l=150000u
+  ad=6.771e+11p pd=3.31e+06u as=0p ps=0u
M1015 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_468_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_129_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_468_264# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_129_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_468_264# C_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1023 VPWR C_N a_468_264# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4_1 A B C D VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=8.7975e+11p ps=6.9e+06u
M1001 a_147_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=3.136e+11p ps=2.8e+06u
M1002 a_345_368# C a_231_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=4.368e+11p ps=3.02e+06u
M1003 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_231_368# B a_147_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y D a_345_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1007 VGND D Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4_2 A B C D VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=9.064e+11p pd=7.51e+06u as=4.44e+11p ps=4.16e+06u
M1001 a_119_368# C a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.216e+11p pd=5.59e+06u as=9.632e+11p ps=8.44e+06u
M1002 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_493_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=7.056e+11p pd=5.74e+06u as=0p ps=0u
M1004 Y D a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1005 Y D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_119_368# D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_493_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1008 a_27_368# C a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_493_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_368# B a_493_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4_4 A B C D VGND VNB VPB VPWR Y
M1000 a_499_368# B a_879_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=1.5568e+12p ps=1.398e+07u
M1001 VGND D Y VNB nlowvt w=740000u l=150000u
+  ad=2.6973e+12p pd=1.469e+07u as=2.4864e+12p ps=1.264e+07u
M1002 Y D a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.608e+11p pd=5.66e+06u as=1.5904e+12p ps=1.404e+07u
M1003 a_27_368# D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_368# D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_879_368# B a_499_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y D a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_499_368# C a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_879_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=8.288e+11p ps=5.96e+06u
M1009 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_499_368# B a_879_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_879_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_368# C a_499_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_879_368# B a_499_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_499_368# C a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_368# C a_499_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_879_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_879_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
M1000 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=8.594e+11p ps=6.85e+06u
M1001 a_347_368# B a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.696e+11p pd=2.9e+06u as=2.688e+11p ps=2.72e+06u
M1002 VGND a_57_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND D_N a_57_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1005 Y a_57_368# a_449_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.48e+11p pd=3.04e+06u as=4.368e+11p ps=3.02e+06u
M1006 a_263_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.06e+11p ps=3.02e+06u
M1007 a_449_368# C a_347_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR D_N a_57_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
M1000 VGND D_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=1.7479e+12p pd=1.217e+07u as=1.824e+11p ps=1.85e+06u
M1001 VPWR D_N a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=5.936e+11p pd=5.36e+06u as=2.8e+11p ps=2.56e+06u
M1002 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=9.879e+11p pd=8.59e+06u as=0p ps=0u
M1003 a_701_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=8.38e+06u as=0p ps=0u
M1004 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_501_368# B a_701_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1006 VGND a_27_392# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_701_368# B a_501_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_701_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_27_392# a_229_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=9.296e+11p ps=8.38e+06u
M1013 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_229_368# a_27_392# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_501_368# C a_229_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_229_368# C a_501_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
M1000 a_781_368# C a_319_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.3496e+12p pd=1.137e+07u as=1.6744e+12p ps=1.419e+07u
M1001 a_319_368# C a_781_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y a_47_88# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.7686e+12p pd=1.662e+07u as=3.0229e+12p ps=2.149e+07u
M1003 VGND a_47_88# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND D_N a_47_88# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.1115e+11p ps=2.85e+06u
M1011 VGND a_47_88# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_47_88# D_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=1.0752e+12p ps=1.004e+07u
M1013 VPWR D_N a_47_88# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_781_368# B a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.5904e+12p ps=1.404e+07u
M1015 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1191_368# B a_781_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_781_368# B a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1191_368# B a_781_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1191_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y a_47_88# a_319_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1023 VPWR A a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y a_47_88# a_319_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_319_368# a_47_88# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_319_368# a_47_88# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_47_88# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_781_368# C a_319_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_319_368# C a_781_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1191_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
M1000 a_611_244# D_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=1.21035e+12p ps=6.39e+06u
M1001 a_400_368# B a_316_368# VPB pshort w=1.12e+06u l=180000u
+  ad=5.432e+11p pd=3.21e+06u as=2.688e+11p ps=2.72e+06u
M1002 a_533_368# a_27_112# a_400_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1003 VGND C_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=1.51135e+12p pd=8.63e+06u as=3.025e+11p ps=2.2e+06u
M1004 a_611_244# D_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1005 Y a_611_244# a_533_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1006 VPWR C_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1007 VGND a_611_244# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.18e+11p ps=4.36e+06u
M1008 Y a_27_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_316_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=2.32715e+12p pd=1.585e+07u as=8.621e+11p ps=8.25e+06u
M1001 Y a_311_124# a_493_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=9.856e+11p ps=8.48e+06u
M1002 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR C_N a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=1.4424e+12p pd=7.06e+06u as=2.8e+11p ps=2.56e+06u
M1004 a_775_368# a_27_392# a_493_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.608e+11p pd=5.66e+06u as=0p ps=0u
M1005 a_493_368# a_27_392# a_775_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_775_368# B a_985_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=9.856e+11p ps=8.48e+06u
M1007 a_493_368# a_311_124# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_985_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_311_124# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_985_368# B a_775_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_27_392# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_985_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_311_124# D_N VGND VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1014 a_311_124# D_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1015 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_311_124# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
M1000 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=1.8722e+12p pd=1.69e+07u as=3.2708e+12p ps=2.364e+07u
M1001 a_119_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.39982e+12p pd=1.162e+07u as=1.8479e+12p ps=1.49e+07u
M1002 a_27_368# B a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_1162_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_1162_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR D_N a_1162_48# VPB pshort w=840000u l=180000u
+  ad=1.5008e+12p pd=1.264e+07u as=2.268e+11p ps=2.22e+06u
M1006 a_1162_48# D_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 a_119_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_864_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_864_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_864_48# C_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1015 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_1162_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR C_N a_864_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_864_48# C_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_900_349# a_864_48# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.6184e+12p pd=1.185e+07u as=0p ps=0u
M1022 a_119_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1162_48# D_N VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_368# a_864_48# a_900_349# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_900_349# a_864_48# a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y a_1162_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_1162_48# a_900_349# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1029 Y a_1162_48# a_900_349# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_900_349# a_1162_48# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_900_349# a_1162_48# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_368# a_864_48# a_900_349# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Y a_864_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_864_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_27_368# B a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_393_74# C1 a_321_74# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=1.554e+11p ps=1.9e+06u
M1001 a_471_74# B1 a_393_74# VNB nlowvt w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=0p ps=0u
M1002 a_82_48# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=6.118e+11p pd=5.03e+06u as=1.20678e+12p ps=8.51e+06u
M1003 VPWR a_82_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1004 VGND A2 a_471_74# VNB nlowvt w=740000u l=150000u
+  ad=4.921e+11p pd=4.29e+06u as=0p ps=0u
M1005 VPWR C1 a_82_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_603_381# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1007 VGND a_82_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.035e+11p ps=2.03e+06u
M1008 a_82_48# D1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_471_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_603_381# A2 a_82_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_321_74# D1 a_82_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.59e+11p ps=2.18e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VPWR D1 a_239_368# VPB pshort w=1e+06u l=180000u
+  ad=1.9396e+12p pd=1.222e+07u as=7.1e+11p ps=5.42e+06u
M1001 VPWR a_239_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1002 a_239_368# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_54_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=7.955e+11p ps=6.59e+06u
M1004 VGND a_239_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 a_461_74# C1 a_369_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=2.294e+11p ps=2.1e+06u
M1006 a_155_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 VGND A1 a_54_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_239_368# D1 a_461_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 X a_239_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_239_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_239_368# A2 a_155_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_239_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_369_74# B1 a_54_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VPWR D1 a_27_392# VPB pshort w=840000u l=180000u
+  ad=2.1934e+12p pd=1.825e+07u as=1.5046e+12p ps=1.239e+07u
M1001 a_287_74# C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=6.6465e+11p ps=6.59e+06u
M1002 a_27_392# A2 a_750_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.9e+11p ps=5.18e+06u
M1003 a_750_392# A2 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_287_74# B1 a_477_198# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.5105e+11p ps=8.36e+06u
M1005 a_477_198# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.295e+12p ps=1.09e+07u
M1006 X a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 a_477_198# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# C1 a_287_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_392# D1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1011 a_27_74# D1 a_27_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B1 a_27_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A1 a_477_198# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_27_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.608e+11p ps=5.66e+06u
M1016 X a_27_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_27_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_750_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_27_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_392# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_27_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A1 a_750_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_392# D1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_392# C1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR C1 a_27_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_477_198# B1 a_287_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_477_198# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_368_74# B1 a_260_74# VNB nlowvt w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=2.886e+11p ps=2.26e+06u
M1001 VPWR A1 a_493_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1872e+12p pd=8.84e+06u as=3.08e+11p ps=2.79e+06u
M1002 VGND A2 a_368_74# VNB nlowvt w=740000u l=150000u
+  ad=3.256e+11p pd=2.36e+06u as=0p ps=0u
M1003 a_493_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.328e+11p ps=5.61e+06u
M1004 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_368_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_182_74# D1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=4.625e+11p ps=2.73e+06u
M1007 a_260_74# C1 a_182_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y D1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_510_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=8.362e+11p pd=8.18e+06u as=4.81e+11p ps=4.26e+06u
M1001 a_40_74# C1 a_299_74# VNB nlowvt w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=5.18e+11p ps=4.36e+06u
M1002 a_299_74# C1 a_40_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A2 a_697_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=9.296e+11p ps=8.38e+06u
M1004 a_510_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_697_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_697_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.6464e+12p pd=1.414e+07u as=0p ps=0u
M1007 a_510_74# B1 a_299_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_697_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_299_74# B1 a_510_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_510_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y D1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR D1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_40_74# D1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1015 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y D1 a_40_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_510_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_954_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=2.8616e+12p pd=1.631e+07u as=2.7776e+12p ps=1.84e+07u
M1001 a_27_74# C1 a_472_74# VNB nlowvt w=740000u l=150000u
+  ad=1.0434e+12p pd=1.022e+07u as=8.288e+11p ps=8.16e+06u
M1002 a_841_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.5688e+12p pd=1.46e+07u as=9.324e+11p ps=8.44e+06u
M1003 a_841_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y D1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.2232e+12p ps=1.517e+07u
M1005 a_841_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_74# C1 a_472_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_472_74# B1 a_841_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_954_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# D1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1011 VGND A1 a_841_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR D1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# D1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_841_74# B1 a_472_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_841_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A2 a_954_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A2 a_841_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A1 a_841_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_472_74# C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_841_74# B1 a_472_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_954_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_472_74# C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A1 a_954_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y D1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A2 a_841_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_954_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_472_74# B1 a_841_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y D1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A2 a_954_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_954_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=2.11e+12p pd=8.4e+06u as=3.136e+11p ps=2.8e+06u
M1001 a_83_264# C1 a_662_136# VNB nlowvt w=640000u l=150000u
+  ad=2.112e+11p pd=1.94e+06u as=2.08e+11p ps=1.93e+06u
M1002 VGND A1 a_257_136# VNB nlowvt w=640000u l=150000u
+  ad=5.891e+11p pd=4.49e+06u as=6.816e+11p ps=4.69e+06u
M1003 a_662_136# B1 a_257_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_401_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1005 a_257_136# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_83_264# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.5e+11p pd=5.1e+06u as=0p ps=0u
M1007 a_83_264# A2 a_401_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B1 a_83_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_195_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=7.498e+11p ps=6.7e+06u
M1001 X a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.4496e+12p ps=9.24e+06u
M1002 VPWR a_27_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 a_195_74# B1 a_117_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1005 a_317_368# A2 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=5.5e+11p ps=5.1e+06u
M1006 a_27_368# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR C1 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_317_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_195_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_117_74# C1 a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR C1 a_91_48# VPB pshort w=840000u l=180000u
+  ad=2.3588e+12p pd=1.71e+07u as=7.736e+11p ps=7.08e+06u
M1001 a_971_391# A2 a_91_48# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1002 VGND a_91_48# X VNB nlowvt w=740000u l=150000u
+  ad=1.1032e+12p pd=1.016e+07u as=4.144e+11p ps=4.08e+06u
M1003 a_91_48# A2 a_971_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_91_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1005 VPWR A1 a_971_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_91_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_91_48# C1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_91_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_91_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_91_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_510_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=8.089e+11p pd=7.65e+06u as=0p ps=0u
M1012 VGND A1 a_510_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_91_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_510_125# B1 a_597_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.032e+11p ps=3.82e+06u
M1015 a_597_125# C1 a_91_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1016 X a_91_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_91_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_971_391# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_597_125# B1 a_510_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_91_48# C1 a_597_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A2 a_510_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_510_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_91_48# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_31_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=2.59e+11p ps=2.18e+06u
M1001 a_311_74# B1 a_31_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1002 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.184e+11p pd=6.12e+06u as=6.72e+11p ps=5.68e+06u
M1003 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1005 Y A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_31_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C1 a_311_74# VNB nlowvt w=740000u l=150000u
+  ad=4.588e+11p pd=2.72e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_303_84# B1 a_30_84# VNB nlowvt w=740000u l=150000u
+  ad=7.067e+11p pd=6.35e+06u as=6.882e+11p ps=6.3e+06u
M1001 a_30_84# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1002 Y C1 a_30_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A2 a_303_84# VNB nlowvt w=740000u l=150000u
+  ad=6.512e+11p pd=6.2e+06u as=0p ps=0u
M1004 a_303_84# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_303_84# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_303_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A2 a_505_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.072e+11p pd=8.34e+06u as=9.296e+11p ps=8.38e+06u
M1008 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.288e+12p ps=1.126e+07u
M1009 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_505_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_505_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_505_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_30_84# B1 a_303_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 a_834_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.0434e+12p ps=1.022e+07u
M1001 Y C1 a_834_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.3664e+12p pd=1.14e+07u as=2.24e+12p ps=1.52e+07u
M1003 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=9.472e+11p pd=8.48e+06u as=1.4578e+12p ps=1.43e+07u
M1004 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_834_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B1 a_834_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_30_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.6464e+12p pd=1.414e+07u as=0p ps=0u
M1012 VPWR A1 a_30_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_30_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_834_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A2 a_30_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_834_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_30_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_834_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_30_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_74# B1 a_834_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A2 a_30_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_30_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_83_244# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=3.13e+11p pd=2.65e+06u as=9.2025e+11p ps=6.03e+06u
M1001 a_320_74# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=3.901e+11p ps=3.89e+06u
M1002 a_320_74# B1 a_83_244# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1003 VPWR a_83_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1004 VPWR A1 a_379_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.9e+11p ps=2.78e+06u
M1005 VGND a_83_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1006 VGND A2 a_320_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_379_387# A2 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VPWR B1 a_247_368# VPB pshort w=1e+06u l=180000u
+  ad=1.204e+12p pd=8.72e+06u as=3.9e+11p ps=2.78e+06u
M1001 a_247_368# A2 a_163_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1002 X a_247_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1003 X a_247_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.14e+11p ps=6.64e+06u
M1004 VPWR a_247_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_54_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=5.032e+11p pd=4.32e+06u as=0p ps=0u
M1006 VGND A1 a_54_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_247_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_163_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_247_368# B1 a_54_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_219_387# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=5.64e+11p pd=4.92e+06u as=1.9384e+12p ps=1.45e+07u
M1001 VGND a_219_387# X VNB nlowvt w=740000u l=150000u
+  ad=1.1573e+12p pd=1.034e+07u as=4.144e+11p ps=4.08e+06u
M1002 X a_219_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=7.744e+11p pd=7.54e+06u as=0p ps=0u
M1004 VGND A2 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_219_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_219_387# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_219_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1008 VPWR B1 a_219_387# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_219_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_125# B1 a_219_387# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1011 a_219_387# A2 a_119_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.4e+11p ps=5.28e+06u
M1012 VPWR a_219_387# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_387# A2 a_219_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A1 a_119_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_119_387# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_219_387# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_219_387# B1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=6.722e+11p ps=3.36e+06u
M1001 a_165_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=7.616e+11p ps=5.84e+06u
M1002 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.32e+11p ps=3.19e+06u
M1003 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1004 Y A2 a_165_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=8.38e+06u as=6.608e+11p ps=5.66e+06u
M1001 a_119_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.608e+11p ps=5.66e+06u
M1002 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.331e+11p pd=2.11e+06u as=8.806e+11p ps=8.3e+06u
M1006 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.069e+11p ps=4.33e+06u
M1008 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=8.399e+11p pd=8.19e+06u as=1.4763e+12p ps=1.435e+07u
M1001 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1003 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.5344e+12p pd=1.394e+07u as=1.3272e+12p ps=1.133e+07u
M1005 VPWR A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.632e+11p pd=8.44e+06u as=0p ps=0u
M1012 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_119_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 X a_203_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=9.926e+11p ps=8.17e+06u
M1001 X a_203_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=5.587e+11p ps=4.44e+06u
M1002 a_119_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1003 a_203_392# A2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=3.9e+11p pd=2.78e+06u as=0p ps=0u
M1004 VPWR a_281_244# a_203_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_203_392# a_281_244# a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=2.176e+11p pd=1.96e+06u as=3.712e+11p ps=3.72e+06u
M1006 VGND B1_N a_281_244# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.75e+11p ps=2.1e+06u
M1007 VPWR B1_N a_281_244# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.982e+11p ps=2.39e+06u
M1008 VGND A1 a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_585_368# A2 a_177_48# VPB pshort w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u
M1001 VGND a_177_48# X VNB nlowvt w=740000u l=150000u
+  ad=7.8915e+11p pd=6.84e+06u as=2.072e+11p ps=2.04e+06u
M1002 VPWR B1_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=1.4348e+12p pd=9.16e+06u as=2.352e+11p ps=2.24e+06u
M1003 VGND A2 a_487_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.07e+11p ps=4.06e+06u
M1004 X a_177_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VPWR a_177_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B1_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5125e+11p ps=1.65e+06u
M1007 X a_177_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_487_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_585_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_177_48# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_487_74# a_27_74# a_177_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.035e+11p ps=2.03e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VPWR A1 a_895_392# VPB pshort w=1e+06u l=180000u
+  ad=2.0896e+12p pd=1.49e+07u as=5.4e+11p ps=5.08e+06u
M1001 X a_193_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1002 VPWR a_193_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_193_48# X VNB nlowvt w=740000u l=150000u
+  ad=1.0914e+12p pd=1.012e+07u as=4.218e+11p ps=4.1e+06u
M1004 VGND A2 a_618_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=7.9445e+11p ps=7.84e+06u
M1005 VGND a_193_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_618_94# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_193_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_193_48# a_27_368# a_618_94# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1009 a_618_94# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1_N a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1011 VPWR a_193_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1 a_618_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_193_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_895_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_618_94# a_27_368# a_193_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_193_48# A2 a_895_392# VPB pshort w=1e+06u l=180000u
+  ad=4.968e+11p pd=4.76e+06u as=0p ps=0u
M1017 a_193_48# a_27_368# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_193_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_27_368# a_193_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND B1_N a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1021 a_895_392# A2 a_193_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR A1 a_398_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.0038e+12p pd=6.52e+06u as=3.36e+11p ps=2.84e+06u
M1001 VGND B1_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=3.6585e+11p pd=3.71e+06u as=1.54e+11p ps=1.66e+06u
M1002 a_308_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.551e+11p pd=4.19e+06u as=0p ps=0u
M1003 a_308_74# a_27_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 VGND A2 a_308_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B1_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 Y a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1007 a_398_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR B1_N a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=1.3578e+12p pd=9.18e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_510_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.104e+11p pd=5.57e+06u as=0p ps=0u
M1002 Y A2 a_510_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1003 a_510_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_225_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=8.88e+11p pd=8.32e+06u as=6.708e+11p ps=6.13e+06u
M1005 a_225_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_225_74# a_27_74# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1008 Y a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_27_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1_N a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1012 VPWR A1 a_510_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_27_74# a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 Y a_828_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=1.6132e+12p ps=1.472e+07u
M1001 a_27_74# a_828_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.3944e+12p pd=1.285e+07u as=1.5904e+12p ps=1.404e+07u
M1003 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.2473e+12p ps=1.099e+07u
M1006 Y a_828_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B1_N a_828_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 Y A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.288e+12p pd=1.126e+07u as=0p ps=0u
M1012 Y a_828_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_828_48# B1_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1014 a_28_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B1_N a_828_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_28_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# a_828_48# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_828_48# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VGND A2 a_245_94# VNB nlowvt w=640000u l=150000u
+  ad=4.931e+11p pd=4.19e+06u as=4.032e+11p ps=3.82e+06u
M1001 a_245_94# B2 a_456_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.576e+11p ps=3.99e+06u
M1002 a_83_264# A2 a_267_392# VPB pshort w=1e+06u l=180000u
+  ad=6.7e+11p pd=5.34e+06u as=2.4e+11p ps=2.48e+06u
M1003 a_245_94# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1005 VPWR B1 a_465_392# VPB pshort w=1e+06u l=180000u
+  ad=1.42e+12p pd=7.02e+06u as=3.9e+11p ps=2.78e+06u
M1006 a_83_264# C1 a_456_74# VNB nlowvt w=640000u l=150000u
+  ad=2.944e+11p pd=2.2e+06u as=0p ps=0u
M1007 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 a_456_74# B1 a_245_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_83_264# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_267_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_465_392# B2 a_83_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VGND a_27_368# X VNB nlowvt w=740000u l=150000u
+  ad=8.325e+11p pd=6.69e+06u as=2.072e+11p ps=2.04e+06u
M1001 a_533_368# A2 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=3.9e+11p pd=2.78e+06u as=6.7e+11p ps=5.34e+06u
M1002 a_27_368# B2 a_335_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1003 a_165_74# B2 a_264_74# VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=4.699e+11p ps=4.23e+06u
M1004 VGND A1 a_264_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A1 a_533_368# VPB pshort w=1e+06u l=180000u
+  ad=1.7732e+12p pd=9.88e+06u as=0p ps=0u
M1006 VPWR C1 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_165_74# C1 a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1008 X a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_264_74# B1 a_165_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_264_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_335_368# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1013 VPWR a_27_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 X a_114_125# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=7.504e+11p pd=5.82e+06u as=2.281e+12p ps=1.709e+07u
M1001 a_27_125# B1 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=7.904e+11p pd=7.59e+06u as=7.456e+11p ps=7.45e+06u
M1002 VGND a_114_125# X VNB nlowvt w=740000u l=150000u
+  ad=1.2421e+12p pd=1.053e+07u as=4.181e+11p ps=4.09e+06u
M1003 X a_114_125# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_300_125# B2 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_114_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_114_125# A2 a_766_387# VPB pshort w=1e+06u l=180000u
+  ad=8.35e+11p pd=7.67e+06u as=6.15e+11p ps=5.23e+06u
M1008 a_300_387# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.85e+11p pd=5.17e+06u as=0p ps=0u
M1009 VGND A2 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_300_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_300_125# B1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_125# C1 a_114_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1013 a_766_387# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_114_125# C1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_114_125# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR C1 a_114_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_766_387# A2 a_114_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_300_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_114_125# B2 a_300_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_114_125# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_300_387# B2 a_114_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_114_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 a_300_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_766_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_125# B2 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_114_125# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_114_125# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 VGND A2 a_239_74# VNB nlowvt w=740000u l=150000u
+  ad=4.736e+11p pd=2.76e+06u as=6.808e+11p ps=6.28e+06u
M1001 a_239_74# B2 a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.217e+11p ps=4.37e+06u
M1002 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.1312e+12p pd=6.5e+06u as=7.504e+11p ps=5.82e+06u
M1003 a_114_74# B1 a_239_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_327_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1005 a_525_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1006 a_239_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B2 a_327_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_525_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_114_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_311_85# B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=1.0841e+12p pd=1.033e+07u as=9.287e+11p ps=8.43e+06u
M1001 a_311_85# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.328e+11p ps=4.4e+06u
M1002 Y B2 a_379_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.24e+11p pd=8.37e+06u as=7e+11p ps=5.73e+06u
M1003 VGND A1 a_311_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# B2 a_311_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A2 a_779_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.608e+11p ps=5.66e+06u
M1006 a_779_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.8032e+12p ps=1.218e+07u
M1007 a_779_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_379_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_379_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_379_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A2 a_311_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_74# B1 a_311_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_779_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_311_85# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1018 a_27_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_311_85# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_27_84# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.4578e+12p pd=1.43e+07u as=4.144e+11p ps=4.08e+06u
M1001 a_1291_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2712e+12p pd=1.123e+07u as=2.5144e+12p ps=2.017e+07u
M1002 a_27_84# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR B1 a_511_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.2656e+12p ps=1.122e+07u
M1004 Y C1 a_27_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_511_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.8984e+12p ps=1.683e+07u
M1006 a_483_74# B2 a_27_84# VNB nlowvt w=740000u l=150000u
+  ad=1.9758e+12p pd=1.866e+07u as=0p ps=0u
M1007 VGND A2 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=9.916e+11p pd=8.6e+06u as=0p ps=0u
M1008 a_483_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_84# B1 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_1291_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_84# B1 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_483_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_483_74# B2 a_27_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_84# B2 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_483_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y C1 a_27_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_511_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A2 a_1291_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_511_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1291_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B2 a_511_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_84# B2 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A1 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR B1 a_511_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A2 a_1291_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_483_74# B1 a_27_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A1 a_483_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_511_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1291_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_483_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y B2 a_511_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_483_74# B1 a_27_84# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1291_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR A1 a_1291_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_299_139# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=5.3175e+11p pd=5.54e+06u as=5.00375e+11p ps=4.3e+06u
M1001 VPWR A1 a_575_392# VPB pshort w=1e+06u l=180000u
+  ad=1.54e+12p pd=7.26e+06u as=3.6e+11p ps=2.72e+06u
M1002 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1003 a_83_260# B1 a_299_139# VNB nlowvt w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=0p ps=0u
M1004 VGND A2 a_299_139# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_401_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1006 a_299_139# B2 a_83_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_83_260# B2 a_401_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1008 a_575_392# A2 a_83_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_578_384# A2 a_82_48# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=3.3e+11p ps=2.66e+06u
M1001 X a_82_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.3128e+12p ps=8.96e+06u
M1002 VPWR a_82_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_82_48# B1 a_307_74# VNB nlowvt w=740000u l=150000u
+  ad=2.294e+11p pd=2.1e+06u as=6.649e+11p ps=6.26e+06u
M1004 X a_82_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=6.5575e+11p ps=6.24e+06u
M1005 VPWR A1 a_578_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_386_384# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1007 a_307_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_82_48# B2 a_386_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_82_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_307_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_307_74# B2 a_82_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VPWR A1 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=2.0354e+12p pd=1.451e+07u as=5.9e+11p ps=5.18e+06u
M1001 a_119_392# A2 a_209_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.4e+11p ps=5.28e+06u
M1002 a_119_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_209_392# A2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_209_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.44e+11p pd=5.63e+06u as=0p ps=0u
M1005 a_27_136# B1 a_209_392# VNB nlowvt w=640000u l=150000u
+  ad=1.0112e+12p pd=9.56e+06u as=3.616e+11p ps=3.69e+06u
M1006 VGND a_209_392# X VNB nlowvt w=740000u l=150000u
+  ad=1.1945e+12p pd=1.055e+07u as=4.144e+11p ps=4.08e+06u
M1007 X a_209_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_209_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_209_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_209_392# B2 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_209_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_136# B2 a_209_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_136# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_209_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_136# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A1 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_209_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_519_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1020 a_209_392# B1 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR B1 a_519_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_519_392# B2 a_209_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_209_392# B2 a_519_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_145_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=2.688e+11p ps=2.72e+06u
M1001 VPWR A1 a_343_368# VPB pshort w=1.12e+06u l=180000u
+  ad=7.616e+11p pd=5.84e+06u as=4.368e+11p ps=3.02e+06u
M1002 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=6.808e+11p ps=6.28e+06u
M1003 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.255e+11p ps=2.63e+06u
M1004 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_145_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_343_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.296e+11p ps=8.38e+06u
M1001 VPWR B1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.608e+11p pd=5.66e+06u as=0p ps=0u
M1002 a_28_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.4282e+12p pd=1.126e+07u as=4.958e+11p ps=4.3e+06u
M1004 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.402e+11p ps=4.42e+06u
M1005 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A2 a_510_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=9.296e+11p ps=8.38e+06u
M1009 a_510_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_510_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_510_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_28_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=2.0566e+12p pd=1.9e+07u as=1.0582e+12p ps=8.78e+06u
M1001 a_120_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=1.7584e+12p ps=1.434e+07u
M1002 a_120_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A1 a_120_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A2 a_120_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2768e+12p pd=1.124e+07u as=0p ps=0u
M1005 a_120_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A2 a_120_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_880_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.3104e+12p pd=1.13e+07u as=0p ps=0u
M1008 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_120_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_880_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=9.768e+11p ps=8.56e+06u
M1012 VPWR A1 a_120_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_880_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B2 a_880_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_880_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_880_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y B2 a_880_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR B1 a_880_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_236_384# A1_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.73e+11p pd=2.33e+06u as=1.6344e+12p ps=9.5e+06u
M1001 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=6.211e+11p pd=4.59e+06u as=2.109e+11p ps=2.05e+06u
M1002 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1003 a_253_94# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1004 a_236_384# A2_N a_253_94# VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1005 a_696_384# B2 a_83_260# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=3.172e+11p ps=2.66e+06u
M1006 a_588_74# a_236_384# a_83_260# VNB nlowvt w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=1.824e+11p ps=1.85e+06u
M1007 a_83_260# a_236_384# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B1 a_696_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_588_74# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A2_N a_236_384# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B2 a_588_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_270_48# A2_N VPWR VPB pshort w=840000u l=180000u
+  ad=3.024e+11p pd=2.4e+06u as=1.68435e+12p ps=1.199e+07u
M1001 X a_204_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=7.087e+11p ps=6.4e+06u
M1002 VPWR A1_N a_270_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_500_74# A2_N a_270_48# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.824e+11p ps=1.85e+06u
M1004 VPWR a_270_48# a_204_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1005 a_204_392# a_270_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=4.699e+11p ps=4.23e+06u
M1006 a_120_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 VGND A1_N a_500_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_204_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 VGND B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_204_392# B2 a_120_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_204_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_204_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR B1 a_41_392# VPB pshort w=1e+06u l=180000u
+  ad=2.2314e+12p pd=1.735e+07u as=8.3e+11p ps=7.66e+06u
M1001 a_41_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_476_48# A2_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1003 VPWR a_313_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=7.224e+11p ps=5.77e+06u
M1004 X a_313_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=1.3531e+12p ps=1.093e+07u
M1005 a_27_74# a_476_48# a_313_392# VNB nlowvt w=640000u l=150000u
+  ad=7.648e+11p pd=7.51e+06u as=2.016e+11p ps=1.91e+06u
M1006 a_313_392# B2 a_41_392# VPB pshort w=1e+06u l=180000u
+  ad=5.556e+11p pd=4.9e+06u as=0p ps=0u
M1007 VPWR A1_N a_476_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_313_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_41_392# B2 a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_476_48# a_313_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_313_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_313_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_313_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_313_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B2 a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A1_N a_835_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1018 VGND a_313_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_313_392# a_476_48# a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_835_94# A2_N a_476_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.952e+11p ps=1.89e+06u
M1021 a_313_392# a_476_48# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B1 a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_74# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_397_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.699e+11p pd=4.23e+06u as=3.896e+11p ps=3.89e+06u
M1001 Y a_134_383# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.30342e+12p ps=8.81e+06u
M1002 VPWR B1 a_493_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1003 a_493_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_134_383# A2_N a_114_74# VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.536e+11p ps=1.76e+06u
M1005 a_134_383# A1_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1006 VPWR A2_N a_134_383# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B2 a_397_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_397_74# a_134_383# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_114_74# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 Y a_136_387# a_518_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.954e+11p ps=8.34e+06u
M1001 a_136_387# A1_N VPWR VPB pshort w=840000u l=180000u
+  ad=5.46225e+11p pd=4.82e+06u as=2.03735e+12p ps=1.491e+07u
M1002 VGND B2 a_518_74# VNB nlowvt w=740000u l=150000u
+  ad=8.869e+11p pd=8.09e+06u as=0p ps=0u
M1003 VPWR A2_N a_136_387# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_799_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1005 Y B2 a_799_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.216e+11p pd=5.59e+06u as=0p ps=0u
M1006 a_518_74# a_136_387# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_134_74# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1008 a_136_387# A2_N a_134_74# VNB nlowvt w=640000u l=150000u
+  ad=2.272e+11p pd=1.99e+06u as=0p ps=0u
M1009 a_799_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_518_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y a_136_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1_N a_134_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B1 a_799_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A1_N a_136_387# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_518_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_136_387# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B1 a_518_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_136_387# A2_N VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_134_74# A2_N a_136_387# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_117_368# A2_N VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=2.7216e+12p ps=2.502e+07u
M1001 Y B2 a_1215_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=1.512e+12p ps=1.39e+07u
M1002 VGND B2 a_857_74# VNB nlowvt w=740000u l=150000u
+  ad=1.3986e+12p pd=1.266e+07u as=1.4578e+12p ps=1.43e+07u
M1003 VPWR A2_N a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1215_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_117_368# A2_N VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_857_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1 a_1215_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A2_N a_117_368# VNB nlowvt w=740000u l=150000u
+  ad=1.1211e+12p pd=1.043e+07u as=4.477e+11p ps=4.17e+06u
M1009 a_857_74# a_117_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1010 VPWR A2_N a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1215_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_74# A1_N VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B1 a_857_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_117_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B1 a_1215_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B1 a_857_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_117_368# A2_N a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_117_368# a_857_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_117_368# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1215_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y a_117_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_368# A2_N a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_857_74# a_117_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_857_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND B2 a_857_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_117_368# A1_N VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A1_N a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_117_368# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_117_368# a_857_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_117_368# A1_N VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y B2 a_1215_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND A1_N a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_74# A1_N VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A1_N a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_857_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR A1_N a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1215_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_857_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_27_74# A2_N a_117_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VGND A1 a_209_74# VNB nlowvt w=640000u l=150000u
+  ad=6.202e+11p pd=4.62e+06u as=8.448e+11p ps=5.2e+06u
M1001 VPWR A1 a_539_387# VPB pshort w=1e+06u l=180000u
+  ad=8.42e+11p pd=5.86e+06u as=3.9e+11p ps=2.78e+06u
M1002 a_209_74# B1 a_131_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1003 a_539_387# A2 a_323_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=9e+11p ps=3.8e+06u
M1004 a_131_74# C1 a_31_387# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1005 a_209_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_31_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VGND A2 a_209_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_31_387# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.5e+11p pd=5.1e+06u as=0p ps=0u
M1009 a_323_387# A3 a_31_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C1 a_31_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_31_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_219_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.958e+11p pd=4.3e+06u as=1.1042e+12p ps=7.58e+06u
M1001 a_135_74# C1 a_32_74# VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=2.701e+11p ps=2.21e+06u
M1002 VGND A3 a_219_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_447_368# A2 a_363_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=2.688e+11p ps=2.72e+06u
M1004 VPWR A1 a_447_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2132e+12p pd=8.73e+06u as=0p ps=0u
M1005 X a_32_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 a_32_74# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=6.736e+11p pd=5.52e+06u as=0p ps=0u
M1007 VPWR C1 a_32_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A1 a_219_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_32_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_363_368# A3 a_32_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_32_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1012 VPWR a_32_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_219_74# B1 a_135_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR C1 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=2.262e+12p pd=1.704e+07u as=1e+12p ps=8e+06u
M1001 X a_83_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=1.5521e+12p ps=1.276e+07u
M1002 VPWR A1 a_1341_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.8e+11p ps=5.36e+06u
M1003 a_83_244# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1341_392# A2 a_1034_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.015e+12p ps=8.03e+06u
M1005 a_1341_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_564_78# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.02922e+12p pd=9.63e+06u as=0p ps=0u
M1007 a_651_78# B1 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=6.88e+11p pd=4.71e+06u as=0p ps=0u
M1008 a_83_244# A3 a_1034_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_83_244# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=8.12e+11p pd=5.93e+06u as=0p ps=0u
M1010 X a_83_244# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_83_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1034_392# A3 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_83_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_83_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_564_78# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1034_392# A2 a_1341_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_83_244# C1 a_651_78# VNB nlowvt w=640000u l=150000u
+  ad=3.4395e+11p pd=2.59e+06u as=0p ps=0u
M1018 VPWR a_83_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_83_244# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B1 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_564_78# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_651_78# C1 a_83_244# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A3 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_83_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_564_78# B1 a_651_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A1 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=7.504e+11p pd=5.82e+06u as=7.504e+11p ps=5.82e+06u
M1001 Y C1 a_469_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.294e+11p ps=2.1e+06u
M1002 a_141_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1003 a_128_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=7.067e+11p ps=4.87e+06u
M1004 a_225_368# A2 a_141_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1005 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_469_74# B1 a_128_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A3 a_225_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_128_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_128_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=9.184e+11p pd=8.36e+06u as=1.232e+12p ps=1.116e+07u
M1001 a_310_368# A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.832e+11p pd=5.7e+06u as=9.744e+11p ps=8.46e+06u
M1002 a_28_368# A2 a_310_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.1174e+12p pd=1.042e+07u as=6.956e+11p ps=6.32e+06u
M1004 a_670_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.18e+11p pd=4.36e+06u as=4.218e+11p ps=4.1e+06u
M1005 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_670_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C1 a_670_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# B1 a_670_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_310_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A3 a_310_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 Y A3 a_841_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.7192e+12p pd=1.203e+07u as=1.7248e+12p ps=1.428e+07u
M1001 VGND A1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=2.19225e+12p pd=1.657e+07u as=1.7316e+12p ps=1.652e+07u
M1002 a_459_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_459_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.02765e+12p ps=1.022e+07u
M1004 VGND A2 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=0p ps=0u
M1006 a_459_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1353_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2656e+12p pd=1.122e+07u as=3.4832e+12p ps=1.966e+07u
M1009 VPWR A1 a_1353_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A3 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A3 a_841_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_459_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1353_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_459_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_74# B1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# B1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_459_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1353_368# A2 a_841_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_841_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_841_368# A2 a_1353_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A3 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_841_368# A2 a_1353_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A2 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1353_368# A2 a_841_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_459_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR A1 a_1353_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_841_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_459_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 a_230_94# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=4.48e+11p pd=3.96e+06u as=6.755e+11p ps=4.76e+06u
M1001 a_84_48# B1 a_230_94# VNB nlowvt w=640000u l=150000u
+  ad=2.272e+11p pd=1.99e+06u as=0p ps=0u
M1002 a_84_48# A3 a_343_368# VPB pshort w=1e+06u l=180000u
+  ad=3.472e+11p pd=2.72e+06u as=3.3e+11p ps=2.66e+06u
M1003 VGND A2 a_230_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_259_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=9.36e+11p ps=5.86e+06u
M1005 VPWR B1 a_84_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_84_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1007 a_230_94# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_84_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_343_368# A2 a_259_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 a_55_264# A3 a_433_392# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=3.9e+11p ps=2.78e+06u
M1001 VPWR B1 a_55_264# VPB pshort w=1e+06u l=180000u
+  ad=1.2386e+12p pd=8.83e+06u as=0p ps=0u
M1002 VGND A2 a_328_74# VNB nlowvt w=740000u l=150000u
+  ad=8.843e+11p pd=6.83e+06u as=6.216e+11p ps=4.64e+06u
M1003 a_55_264# B1 a_328_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1004 X a_55_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.64e+11p pd=2.89e+06u as=0p ps=0u
M1005 VGND a_55_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1006 X a_55_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_349_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1008 a_328_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_433_392# A2 a_349_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_328_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_55_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_971_392# VPB pshort w=1e+06u l=180000u
+  ad=1.6046e+12p pd=1.373e+07u as=5.8e+11p ps=5.16e+06u
M1001 a_971_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_86_260# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1003 VGND a_86_260# X VNB nlowvt w=740000u l=150000u
+  ad=1.2225e+12p pd=1.183e+07u as=4.144e+11p ps=4.08e+06u
M1004 VPWR B1 a_86_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_699_392# A2 a_971_392# VPB pshort w=1e+06u l=180000u
+  ad=8.4e+11p pd=7.68e+06u as=0p ps=0u
M1006 X a_86_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_86_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.048e+11p ps=5.56e+06u
M1008 X a_86_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_492_125# B1 a_86_260# VNB nlowvt w=640000u l=150000u
+  ad=1.0624e+12p pd=9.72e+06u as=2.112e+11p ps=1.94e+06u
M1010 VGND A2 a_492_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_86_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_86_260# A3 a_699_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_699_392# A3 a_86_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_86_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_971_392# A2 a_699_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_492_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_492_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_86_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_492_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_86_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A3 a_492_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_492_125# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_86_260# B1 a_492_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_206_368# A2 a_122_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=2.688e+11p ps=2.72e+06u
M1001 a_114_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.292e+11p pd=4.12e+06u as=9.093e+11p ps=5.45e+06u
M1002 Y B1 a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=2.479e+11p pd=2.15e+06u as=0p ps=0u
M1003 a_122_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.272e+11p ps=5.6e+06u
M1004 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=7.392e+11p ps=3.56e+06u
M1005 a_114_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A3 a_206_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.296e+11p ps=8.38e+06u
M1001 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_300_368# A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1003 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=1.2616e+12p pd=7.93e+06u as=1.0582e+12p ps=1.026e+07u
M1004 a_28_368# A2 a_300_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=0p ps=0u
M1008 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_300_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=9.856e+11p ps=8.48e+06u
M1010 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A3 a_300_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VGND A1 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=2.2892e+12p pd=1.54e+07u as=1.924e+12p ps=1.852e+07u
M1001 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.7976e+12p pd=9.93e+06u as=1.8928e+12p ps=1.458e+07u
M1002 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A2 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_82# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A1 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_490_368# A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2656e+12p pd=1.122e+07u as=0p ps=0u
M1009 a_28_368# A2 a_490_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_82# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_82# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.288e+12p pd=1.126e+07u as=0p ps=0u
M1013 Y B1 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1014 VGND A3 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y B1 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_490_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_82# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A3 a_27_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_490_368# A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_82# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A3 a_490_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_28_368# A2 a_490_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_82# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_490_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_82# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_82# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A3 a_490_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_251_74# B1 a_83_264# VNB nlowvt w=640000u l=150000u
+  ad=6.176e+11p pd=5.77e+06u as=2.848e+11p ps=2.17e+06u
M1001 a_551_368# B2 a_83_264# VPB pshort w=1e+06u l=180000u
+  ad=4.15e+11p pd=2.83e+06u as=3.6e+11p ps=2.72e+06u
M1002 VGND A2 a_251_74# VNB nlowvt w=640000u l=150000u
+  ad=5.626e+11p pd=4.44e+06u as=0p ps=0u
M1003 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=7.996e+11p pd=5.76e+06u as=3.136e+11p ps=2.8e+06u
M1004 VPWR B1 a_551_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_251_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1006 a_83_264# B2 a_251_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1008 a_251_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_335_368# A2 a_251_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=0p ps=0u
M1010 a_251_74# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_83_264# A3 a_335_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_433_368# A2 a_349_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=2.4e+11p ps=2.48e+06u
M1001 a_83_264# B2 a_349_74# VNB nlowvt w=740000u l=150000u
+  ad=6.771e+11p pd=3.31e+06u as=7.289e+11p ps=6.41e+06u
M1002 a_349_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=9.62e+11p ps=7.04e+06u
M1003 a_655_368# B2 a_83_264# VPB pshort w=1e+06u l=180000u
+  ad=3.9e+11p pd=2.78e+06u as=3.9e+11p ps=2.78e+06u
M1004 X a_83_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1436e+12p ps=8.64e+06u
M1005 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_83_264# A3 a_433_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_349_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B1 a_655_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_349_74# B1 a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1011 VGND A2 a_349_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_349_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_961_392# A3 a_83_256# VPB pshort w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.6e+11p ps=5.12e+06u
M1001 a_1237_392# A2 a_961_392# VPB pshort w=1e+06u l=180000u
+  ad=7.3e+11p pd=5.46e+06u as=0p ps=0u
M1002 a_564_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.2032e+12p pd=1.144e+07u as=1.5408e+12p ps=1.279e+07u
M1003 VPWR a_83_256# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.7126e+12p pd=1.394e+07u as=7.392e+11p ps=5.8e+06u
M1004 a_564_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A1 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_83_256# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_256# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_83_256# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_83_256# B1 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=0p ps=0u
M1011 a_1237_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A3 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_961_392# A2 a_1237_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_564_74# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_83_256# VGND VNB nlowvt w=740000u l=150000u
+  ad=5.069e+11p pd=4.33e+06u as=0p ps=0u
M1016 a_83_256# B2 a_537_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.8e+11p ps=5.36e+06u
M1017 a_83_256# A3 a_961_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_537_388# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_537_388# B2 a_83_256# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_83_256# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_564_74# B2 a_83_256# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_83_256# B2 a_564_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 a_537_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_83_256# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_564_74# B1 a_83_256# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A1 a_1237_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_83_256# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=5.439e+11p pd=4.43e+06u as=6.771e+11p ps=6.27e+06u
M1001 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_345_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=5.264e+11p ps=3.18e+06u
M1003 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=2.65e+06u
M1004 VPWR A1 a_459_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.72e+11p pd=5.68e+06u as=4.368e+11p ps=3.02e+06u
M1005 a_459_368# A2 a_345_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_131_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1007 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B2 a_131_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 a_771_368# A2 a_499_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.104e+11p pd=5.57e+06u as=9.296e+11p ps=8.38e+06u
M1001 a_499_368# A2 a_771_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.296e+11p ps=8.38e+06u
M1003 a_27_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.856e+11p pd=8.48e+06u as=0p ps=0u
M1005 a_27_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_771_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.4208e+12p pd=1.272e+07u as=1.5162e+12p ps=8.64e+06u
M1008 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_771_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1012 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A3 a_499_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_499_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=2.9524e+12p pd=2.427e+07u as=9.435e+11p ps=8.47e+06u
M1001 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.7051e+12p ps=1.361e+07u
M1002 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_1333_368# A2 a_861_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2656e+12p pd=1.122e+07u as=1.7584e+12p ps=1.434e+07u
M1004 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A3 a_861_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2096e+12p pd=1.112e+07u as=0p ps=0u
M1007 a_861_368# A2 a_1333_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_861_368# A2 a_1333_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1333_368# A2 a_861_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.5344e+12p pd=1.394e+07u as=1.6576e+12p ps=1.416e+07u
M1013 a_861_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_368# B2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1333_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1333_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A1 a_1333_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A3 a_861_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y B2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A1 a_1333_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_861_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR a_83_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.3554e+12p pd=7.11e+06u as=3.136e+11p ps=2.8e+06u
M1001 VGND A4 a_326_74# VNB nlowvt w=640000u l=150000u
+  ad=8.899e+11p pd=6.71e+06u as=6.24e+11p ps=5.79e+06u
M1002 a_83_270# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=3.7225e+11p pd=2.95e+06u as=0p ps=0u
M1003 a_446_368# A4 a_83_270# VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1004 a_326_74# B1 a_83_270# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1005 a_644_368# A2 a_530_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=4.368e+11p ps=3.02e+06u
M1006 VGND A2 a_326_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_530_368# A3 a_446_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_326_74# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_644_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_83_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 a_326_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_27_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=6.364e+11p pd=6.16e+06u as=1.2691e+12p ps=9.35e+06u
M1001 X a_431_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1002 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=1.6872e+12p ps=9.9e+06u
M1003 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR B1 a_431_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.236e+11p ps=3.02e+06u
M1005 a_203_368# A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1006 a_431_368# A4 a_317_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.368e+11p ps=3.02e+06u
M1007 VGND a_431_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_317_368# A3 a_203_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_431_368# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1010 X a_431_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1011 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_431_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_523_124# A4 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.1456e+12p pd=1.126e+07u as=1.69995e+12p ps=1.463e+07u
M1001 a_1216_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.608e+11p pd=5.66e+06u as=1.5693e+12p ps=1.363e+07u
M1002 a_762_368# A2 a_1216_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.856e+11p pd=8.48e+06u as=0p ps=0u
M1003 X a_110_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1004 a_523_124# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_523_124# B1 a_110_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 VPWR a_110_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_110_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_523_124# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_110_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_110_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1011 a_110_48# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=5.404e+11p pd=5.02e+06u as=0p ps=0u
M1012 a_523_124# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B1 a_110_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_854_368# A3 a_762_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1016 a_110_48# B1 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_110_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A3 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_110_48# A4 a_854_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_110_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_854_368# A4 a_110_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_762_368# A3 a_854_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_110_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1216_368# A2 a_762_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A1 a_1216_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A4 a_523_124# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_157_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=7.104e+11p pd=6.36e+06u as=6.327e+11p ps=4.67e+06u
M1001 a_475_368# A2 a_361_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=4.368e+11p ps=3.02e+06u
M1002 a_361_368# A3 a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.472e+11p ps=2.86e+06u
M1003 a_157_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_475_368# VPB pshort w=1.12e+06u l=180000u
+  ad=8.736e+11p pd=6.04e+06u as=0p ps=0u
M1005 a_263_368# A4 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=2.88e+06u
M1006 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_157_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A4 a_157_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_157_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_314_368# A3 a_610_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.0472e+12p pd=8.59e+06u as=6.048e+11p ps=5.56e+06u
M1001 VPWR A1 a_807_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.016e+11p pd=8.33e+06u as=9.072e+11p ps=8.34e+06u
M1002 a_132_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.4245e+12p pd=1.273e+07u as=1.0397e+12p ps=8.73e+06u
M1003 a_807_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A4 a_132_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_132_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1006 VGND A3 a_132_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_132_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A4 a_314_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1009 a_132_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_314_368# A4 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_132_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_610_368# A2 a_807_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1 a_132_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_807_368# A2 a_610_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A2 a_132_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B1 a_132_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_610_368# A3 a_314_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 VGND A4 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.1756e+12p pd=1.772e+07u as=2.3976e+12p ps=2.276e+07u
M1001 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_339_368# A3 a_791_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.5344e+12p pd=1.394e+07u as=1.3216e+12p ps=1.132e+07u
M1004 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.344e+12p pd=1.136e+07u as=1.0192e+12p ps=8.54e+06u
M1005 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A4 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1010 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_791_368# A2 a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=1.5344e+12p ps=1.394e+07u
M1014 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A4 a_339_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1191_368# A2 a_791_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_339_368# A4 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_791_368# A2 a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A4 a_339_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_339_368# A3 a_791_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1191_368# A2 a_791_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_339_368# A4 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_791_368# A3 a_339_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A1 a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1191_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_791_368# A3 a_339_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A1 a_1191_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1191_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2_1 A B VGND VNB VPB VPWR X
M1000 X a_63_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=5.7345e+11p ps=4.42e+06u
M1001 a_155_368# B a_63_368# VPB pshort w=840000u l=180000u
+  ad=2.016e+11p pd=2.16e+06u as=2.352e+11p ps=2.24e+06u
M1002 VGND A a_63_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.6125e+11p ps=2.05e+06u
M1003 a_63_368# B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_63_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=6.398e+11p ps=3.46e+06u
M1005 VPWR A a_155_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2_2 A B VGND VNB VPB VPWR X
M1000 VPWR A a_117_368# VPB pshort w=1e+06u l=180000u
+  ad=7.072e+11p pd=5.76e+06u as=2.1e+11p ps=2.42e+06u
M1001 VGND a_27_368# X VNB nlowvt w=740000u l=150000u
+  ad=6.823e+11p pd=6.18e+06u as=2.072e+11p ps=2.04e+06u
M1002 X a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.248e+11p pd=2.82e+06u as=0p ps=0u
M1003 a_27_368# B VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1004 a_117_368# B a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 VGND A a_27_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_27_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2_4 A B VGND VNB VPB VPWR X
M1000 VGND B a_83_260# VNB nlowvt w=740000u l=150000u
+  ad=1.6058e+12p pd=1.026e+07u as=2.479e+11p ps=2.15e+06u
M1001 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.3096e+12p ps=1.114e+07u
M1002 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_83_260# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_496_388# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1006 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_83_260# B a_496_388# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1008 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=0p ps=0u
M1009 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_496_388# B a_83_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A a_496_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2b_1 A B_N VGND VNB VPB VPWR X
M1000 a_264_368# a_27_112# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=7.357e+11p ps=5.01e+06u
M1001 VGND A a_264_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_264_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=7.218e+11p ps=5.39e+06u
M1003 VGND B_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=3.685e+11p ps=2.44e+06u
M1004 a_356_368# a_27_112# a_264_368# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1005 VPWR B_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 VPWR A a_356_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_264_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2b_2 A B_N VGND VNB VPB VPWR X
M1000 a_187_48# a_27_368# a_473_368# VPB pshort w=1e+06u l=180000u
+  ad=4e+11p pd=2.8e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR B_N a_27_368# VPB pshort w=840000u l=180000u
+  ad=8.002e+11p pd=5.97e+06u as=2.352e+11p ps=2.24e+06u
M1002 VGND B_N a_27_368# VNB nlowvt w=550000u l=150000u
+  ad=9.5555e+11p pd=7.08e+06u as=1.5675e+11p ps=1.67e+06u
M1003 a_187_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=2.208e+11p pd=1.97e+06u as=0p ps=0u
M1004 X a_187_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VGND a_187_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_473_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_27_368# a_187_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_187_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.432e+11p ps=3.21e+06u
M1009 X a_187_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2b_4 A B_N VGND VNB VPB VPWR X
M1000 a_81_296# A VGND VNB nlowvt w=640000u l=150000u
+  ad=4.672e+11p pd=4.02e+06u as=1.1509e+12p ps=1.032e+07u
M1001 a_81_296# a_676_48# a_492_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=8.2e+11p ps=7.64e+06u
M1002 a_492_392# a_676_48# a_81_296# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_492_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.5272e+12p ps=1.358e+07u
M1004 VPWR A a_492_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_81_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=4.13e+06u
M1006 a_81_296# a_676_48# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_81_296# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_81_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1009 VPWR a_81_296# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_81_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_81_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_81_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_81_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_676_48# B_N VGND VNB nlowvt w=640000u l=150000u
+  ad=6.272e+11p pd=3.24e+06u as=0p ps=0u
M1015 a_676_48# B_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1016 VPWR a_81_296# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_676_48# a_81_296# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or3_1 A B C VGND VNB VPB VPWR X
M1000 a_119_368# C a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1001 VGND A a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=4.71e+11p pd=4.12e+06u as=5.225e+11p ps=4.1e+06u
M1002 a_203_368# B a_119_368# VPB pshort w=1e+06u l=180000u
+  ad=3.9e+11p pd=2.78e+06u as=0p ps=0u
M1003 a_27_74# B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=7.3e+11p ps=3.64e+06u
M1005 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 VPWR A a_203_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or3_2 A B C VGND VNB VPB VPWR X
M1000 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=9.725e+11p pd=7.09e+06u as=2.072e+11p ps=2.04e+06u
M1001 VPWR A a_237_392# VPB pshort w=1e+06u l=180000u
+  ad=8.296e+11p pd=6e+06u as=3.9e+11p ps=2.78e+06u
M1002 a_237_392# B a_153_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1003 a_153_392# C a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1004 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VGND A a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.064e+11p ps=3.83e+06u
M1006 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or3_4 A B C VGND VNB VPB VPWR X
M1000 X a_305_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=9.879e+11p ps=8.59e+06u
M1001 VGND A a_305_388# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.625e+11p ps=4.21e+06u
M1002 VGND a_305_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_305_388# C a_209_388# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=6.25e+11p ps=5.25e+06u
M1004 X a_305_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.2816e+12p ps=1.109e+07u
M1005 a_209_388# C a_305_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_119_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.9e+11p ps=5.18e+06u
M1007 VPWR a_305_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C a_305_388# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_388# B a_209_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_305_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_305_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_305_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_388# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_209_388# B a_119_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_305_388# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_305_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or3b_1 A B C_N VGND VNB VPB VPWR X
M1000 a_239_74# B VGND VNB nlowvt w=550000u l=150000u
+  ad=3.3e+11p pd=3.4e+06u as=8.0375e+11p ps=6.43e+06u
M1001 a_455_391# B a_371_391# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.4e+11p ps=2.48e+06u
M1002 VGND A a_239_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_239_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=7.134e+11p ps=5.37e+06u
M1004 VGND a_127_74# a_239_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_455_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_239_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 a_127_74# C_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.595e+11p pd=1.68e+06u as=0p ps=0u
M1008 a_127_74# C_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.436e+11p pd=2.26e+06u as=0p ps=0u
M1009 a_371_391# a_127_74# a_239_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or3b_2 A B C_N VGND VNB VPB VPWR X
M1000 a_190_260# a_27_368# VGND VNB nlowvt w=640000u l=150000u
+  ad=4.064e+11p pd=3.83e+06u as=9.1395e+11p ps=6.95e+06u
M1001 a_461_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=9.8195e+11p ps=6.3e+06u
M1002 VPWR C_N a_27_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1003 a_545_368# B a_461_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=0p ps=0u
M1004 X a_190_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VGND C_N a_27_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1006 VGND B a_190_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_190_260# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_190_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_190_260# a_27_368# a_545_368# VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1010 X a_190_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1011 VPWR a_190_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or3b_4 A B C_N VGND VNB VPB VPWR X
M1000 VPWR A a_220_392# VPB pshort w=1e+06u l=180000u
+  ad=1.2948e+12p pd=1.112e+07u as=6e+11p ps=5.2e+06u
M1001 X a_412_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.329e+11p pd=4.13e+06u as=1.64125e+12p ps=1.215e+07u
M1002 X a_412_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_412_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.048e+11p ps=5.56e+06u
M1004 a_412_392# a_27_392# a_310_392# VPB pshort w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=6e+11p ps=5.2e+06u
M1005 VPWR C_N a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1006 a_412_392# B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 VGND a_412_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_310_392# a_27_392# a_412_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_392# a_412_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_220_392# B a_310_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_220_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A a_412_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_310_392# B a_220_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_412_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND C_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1016 VPWR a_412_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_412_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_412_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4_1 A B C D VGND VNB VPB VPWR X
M1000 X a_44_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=5.4e+11p ps=3.26e+06u
M1001 a_136_392# D a_44_392# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1002 VGND C a_44_392# VNB nlowvt w=550000u l=150000u
+  ad=7.822e+11p pd=6.34e+06u as=3.96e+11p ps=3.64e+06u
M1003 a_44_392# D VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_44_392# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_334_392# B a_220_392# VPB pshort w=1e+06u l=180000u
+  ad=3.9e+11p pd=2.78e+06u as=3.9e+11p ps=2.78e+06u
M1006 a_44_392# B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_44_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 a_220_392# C a_136_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_334_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4_2 A B C D VGND VNB VPB VPWR X
M1000 a_261_392# C a_177_392# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.4e+11p ps=2.48e+06u
M1001 a_345_392# B a_261_392# VPB pshort w=1e+06u l=180000u
+  ad=4e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_85_392# B VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=1.24458e+12p ps=9.28e+06u
M1003 X a_85_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 a_85_392# D VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A a_85_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C a_85_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_85_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_85_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=8.142e+11p ps=5.95e+06u
M1009 VPWR a_85_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_177_392# D a_85_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1011 VPWR A a_345_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4_4 A B C D VGND VNB VPB VPWR X
M1000 a_83_264# D a_965_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=5.9e+11p ps=5.18e+06u
M1001 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=2.2402e+12p pd=1.413e+07u as=6.549e+11p ps=4.73e+06u
M1002 a_965_392# D a_83_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_499_392# C a_965_392# VPB pshort w=1e+06u l=180000u
+  ad=9.3e+11p pd=7.86e+06u as=0p ps=0u
M1004 a_83_264# B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1005 X a_83_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.1996e+12p ps=1.092e+07u
M1006 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_591_392# B a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1015 a_83_264# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_591_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_591_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_499_392# B a_591_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_965_392# C a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4b_1 A B C D_N VGND VNB VPB VPWR X
M1000 VGND C a_228_74# VNB nlowvt w=550000u l=150000u
+  ad=7.8175e+11p pd=6.35e+06u as=6.6275e+11p ps=4.61e+06u
M1001 VPWR D_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=8.268e+11p pd=5.6e+06u as=2.352e+11p ps=2.24e+06u
M1002 X a_228_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 a_527_368# B a_443_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=2.4e+11p ps=2.48e+06u
M1004 VPWR A a_527_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_228_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1006 a_228_74# B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_359_368# a_27_74# a_228_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1008 VGND D_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 a_443_368# C a_359_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_228_74# a_27_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A a_228_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4b_2 A B C D_N VGND VNB VPB VPWR X
M1000 a_455_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=9.216e+11p ps=6.22e+06u
M1001 a_641_392# C a_539_392# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=3.3e+11p ps=2.66e+06u
M1002 a_190_48# C VGND VNB nlowvt w=640000u l=150000u
+  ad=4.896e+11p pd=4.09e+06u as=1.10645e+12p ps=8.83e+06u
M1003 VPWR D_N a_27_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1004 a_190_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_190_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 a_190_48# a_27_368# a_641_392# VPB pshort w=1e+06u l=180000u
+  ad=4.3e+11p pd=2.86e+06u as=0p ps=0u
M1007 a_539_392# B a_455_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B a_190_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_190_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1010 VGND D_N a_27_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1011 VGND a_27_368# a_190_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_190_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_190_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4b_4 A B C D_N VGND VNB VPB VPWR X
M1000 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=1.3615e+12p pd=1.11e+07u as=5.069e+11p ps=4.33e+06u
M1001 a_119_392# B a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=8.8e+11p ps=7.76e+06u
M1002 VPWR A a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=1.269e+12p pd=1.106e+07u as=0p ps=0u
M1003 a_499_392# C a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1004 a_27_74# a_563_48# a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 a_27_392# B a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_119_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_499_392# a_563_48# a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_392# C a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND D_N a_563_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.2135e+11p ps=2.98e+06u
M1012 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.2395e+12p ps=7.79e+06u
M1014 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1015 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# a_563_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR D_N a_563_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1020 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
M1000 a_357_378# a_219_424# VGND VNB nlowvt w=550000u l=150000u
+  ad=3.7675e+11p pd=3.57e+06u as=9.22e+11p ps=7.96e+06u
M1001 a_629_378# B a_533_378# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=3e+11p ps=2.6e+06u
M1002 a_533_378# a_27_424# a_449_378# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1003 a_219_424# D_N VPWR VPB pshort w=840000u l=180000u
+  ad=4.2525e+11p pd=2.94e+06u as=7.094e+11p ps=5.37e+06u
M1004 VGND C_N a_27_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1005 VPWR C_N a_27_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 VPWR A a_629_378# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_357_378# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1008 a_219_424# D_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1009 VGND A a_357_378# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_357_378# B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_357_378# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_449_378# a_219_424# a_357_378# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1013 VGND a_27_424# a_357_378# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
M1000 VGND a_548_110# a_182_270# VNB nlowvt w=640000u l=150000u
+  ad=1.16472e+12p pd=9.37e+06u as=5.192e+11p ps=4.27e+06u
M1001 VPWR A a_692_392# VPB pshort w=1e+06u l=180000u
+  ad=9.926e+11p pd=8.39e+06u as=2.1e+11p ps=2.42e+06u
M1002 a_692_392# B a_590_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1003 a_182_270# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_548_110# C_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.31e+11p pd=2.23e+06u as=0p ps=0u
M1005 X a_182_270# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 X a_182_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1007 VGND a_182_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND D_N a_27_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 VPWR a_182_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_548_110# C_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1011 a_506_392# a_27_424# a_182_270# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.7e+11p ps=2.54e+06u
M1012 a_590_392# a_548_110# a_506_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A a_182_270# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_182_270# a_27_424# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR D_N a_27_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
M1000 a_1273_392# B a_1063_392# VPB pshort w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.9e+11p ps=5.18e+06u
M1001 VGND a_193_277# X VNB nlowvt w=740000u l=150000u
+  ad=2.0924e+12p pd=1.558e+07u as=6.919e+11p ps=4.83e+06u
M1002 a_1273_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.5228e+12p ps=1.154e+07u
M1003 X a_193_277# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.184e+11p pd=6.12e+06u as=0p ps=0u
M1004 VPWR A a_1273_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_193_277# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_193_277# a_27_94# a_791_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=8.3e+11p ps=7.66e+06u
M1007 VGND A a_193_277# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.4134e+12p ps=6.78e+06u
M1008 VGND D_N a_27_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1009 a_681_368# C_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.719e+11p pd=1.85e+06u as=0p ps=0u
M1010 a_791_392# a_27_94# a_193_277# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR D_N a_27_94# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1012 X a_193_277# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_193_277# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_193_277# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_193_277# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_791_392# a_681_368# a_1063_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_193_277# a_27_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1063_392# a_681_368# a_791_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_193_277# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_193_277# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_681_368# a_193_277# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_681_368# C_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1023 a_1063_392# B a_1273_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 a_353_93# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=2.8826e+12p ps=2.42e+07u
M1001 a_1906_424# a_977_243# VPWR VPB pshort w=840000u l=180000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1002 a_305_119# D a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.129e+11p ps=3.17e+06u
M1003 a_197_119# a_867_82# a_1162_497# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1004 VGND RESET_B a_1579_258# VNB nlowvt w=420000u l=150000u
+  ad=2.11888e+12p pd=1.742e+07u as=1.197e+11p ps=1.41e+06u
M1005 a_977_243# a_1162_497# a_1434_78# VNB nlowvt w=550000u l=150000u
+  ad=2.09e+11p pd=1.86e+06u as=5.1045e+11p ps=4.25e+06u
M1006 a_119_119# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 Q_N a_2133_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 VPWR SCD a_27_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=3.552e+11p ps=3.67e+06u
M1009 a_2392_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.947e+11p pd=4.37e+06u as=0p ps=0u
M1010 VGND a_2133_410# a_2164_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1011 a_197_119# D a_215_464# VPB pshort w=640000u l=180000u
+  ad=3.84e+11p pd=3.76e+06u as=1.536e+11p ps=1.76e+06u
M1012 VPWR a_2133_410# a_2091_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 a_27_464# a_353_93# a_197_119# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1162_497# a_867_82# a_1084_497# VPB pshort w=420000u l=180000u
+  ad=2.107e+11p pd=1.99e+06u as=8.82e+10p ps=1.26e+06u
M1015 a_1954_119# a_867_82# a_1906_424# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=0p ps=0u
M1016 VPWR a_2133_410# a_3078_384# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1017 a_197_119# a_662_82# a_1162_497# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND CLK_N a_662_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1019 a_867_82# a_662_82# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.219e+11p pd=2.35e+06u as=0p ps=0u
M1020 a_1162_497# a_662_82# a_1151_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1021 a_353_93# SCE VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1022 Q a_3078_384# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1023 a_2512_392# a_1579_258# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1024 VGND a_2133_410# a_3078_384# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1025 a_1151_119# a_977_243# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND SET_B a_1434_78# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1954_119# a_662_82# a_1876_119# VNB nlowvt w=550000u l=150000u
+  ad=4.807e+11p pd=2.9e+06u as=1.32e+11p ps=1.58e+06u
M1028 VPWR SET_B a_2133_410# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1029 VPWR CLK_N a_662_82# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1030 a_2091_508# a_662_82# a_1954_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1084_497# a_977_243# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2392_74# a_1954_119# a_2133_410# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.812e+11p ps=2.24e+06u
M1033 a_867_82# a_662_82# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1034 a_197_119# SCE a_119_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_353_93# a_305_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_215_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1531_424# a_1162_497# a_977_243# VPB pshort w=840000u l=180000u
+  ad=2.016e+11p pd=2.16e+06u as=6.09e+11p ps=4.81e+06u
M1038 Q a_3078_384# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1039 a_2133_410# a_1579_258# a_2392_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_2164_119# a_867_82# a_1954_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_1579_258# a_1531_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1876_119# a_977_243# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Q_N a_2133_410# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1044 a_977_243# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1434_78# a_1579_258# a_977_243# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_2133_410# a_1954_119# a_2512_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR RESET_B a_1579_258# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=3.529e+11p ps=3.68e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 VPWR RESET_B a_1643_257# VPB pshort w=640000u l=180000u
+  ad=3.89413e+12p pd=2.968e+07u as=1.792e+11p ps=1.84e+06u
M1001 a_871_368# a_688_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_2174_508# a_688_98# a_1997_82# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=2.667e+11p ps=2.39e+06u
M1003 a_1157_464# a_871_368# a_1073_464# VPB pshort w=420000u l=180000u
+  ad=2.107e+11p pd=1.99e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_1595_424# a_1157_464# a_1007_366# VPB pshort w=840000u l=180000u
+  ad=2.016e+11p pd=2.16e+06u as=9.702e+11p ps=5.67e+06u
M1005 VPWR SET_B a_2216_410# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1006 a_2452_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=5.7435e+11p pd=4.64e+06u as=2.86405e+12p ps=2.37e+07u
M1007 VGND a_2216_410# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1008 a_119_119# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 a_197_119# a_871_368# a_1157_464# VNB nlowvt w=420000u l=150000u
+  ad=4.347e+11p pd=3.75e+06u as=1.281e+11p ps=1.45e+06u
M1010 VGND RESET_B a_1643_257# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1011 a_2452_74# a_1997_82# a_2216_410# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1012 VPWR SCD a_27_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1013 a_209_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1014 VPWR a_2216_410# a_3272_94# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1015 a_2247_82# a_871_368# a_1997_82# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=4.945e+11p ps=3.3e+06u
M1016 a_1157_464# a_688_98# a_1185_125# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 a_341_410# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1018 a_197_119# a_688_98# a_1157_464# VPB pshort w=640000u l=180000u
+  ad=3.84e+11p pd=3.76e+06u as=0p ps=0u
M1019 a_1007_366# a_1157_464# a_1473_73# VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=6.0335e+11p ps=4.55e+06u
M1020 a_1473_73# a_1643_257# a_1007_366# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_2216_410# a_3272_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1022 a_1989_424# a_1007_366# VPWR VPB pshort w=840000u l=180000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1023 a_1997_82# a_688_98# a_1902_125# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.16375e+11p ps=2.18e+06u
M1024 Q_N a_2216_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_3272_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1026 Q_N a_2216_410# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 a_1997_82# a_871_368# a_1989_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_341_410# a_363_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1029 Q a_3272_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1030 a_1073_464# a_1007_366# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1185_125# a_1007_366# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_2216_410# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1643_257# a_1595_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2559_392# a_1643_257# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1035 VPWR a_3272_94# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_2216_410# a_2174_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_197_119# SCE a_119_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND CLK_N a_688_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1039 a_341_410# SCE VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1040 a_2216_410# a_1997_82# a_2559_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_2216_410# a_1643_257# a_2452_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_197_119# D a_209_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND a_3272_94# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_363_119# D a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_27_464# a_341_410# a_197_119# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_871_368# a_688_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1047 VGND a_2216_410# a_2247_82# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VPWR CLK_N a_688_98# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1049 a_1902_125# a_1007_366# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_1007_366# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VGND SET_B a_1473_73# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q
+ Q_N
M1000 VGND a_1250_231# a_1192_96# VNB nlowvt w=420000u l=150000u
+  ad=2.22013e+12p pd=1.787e+07u as=1.61875e+11p ps=1.78e+06u
M1001 VGND a_2037_442# a_2061_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1002 a_877_98# a_622_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1003 a_1881_420# a_877_98# a_1880_119# VNB nlowvt w=550000u l=150000u
+  ad=2.3445e+11p pd=2.34e+06u as=1.155e+11p ps=1.52e+06u
M1004 a_2271_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=0p ps=0u
M1005 Q a_2881_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 a_119_119# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 VGND RESET_B a_1625_93# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1008 VPWR a_1625_93# a_1583_379# VPB pshort w=840000u l=180000u
+  ad=2.88865e+12p pd=2.393e+07u as=2.016e+11p ps=2.16e+06u
M1009 VPWR a_1625_93# a_2387_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1010 VPWR SCD a_27_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1011 a_299_119# D a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.709e+11p ps=2.97e+06u
M1012 a_1881_420# a_622_98# a_1769_379# VPB pshort w=840000u l=180000u
+  ad=2.709e+11p pd=2.4e+06u as=3.438e+11p ps=2.85e+06u
M1013 Q_N a_2037_442# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1014 VPWR CLK a_622_98# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1015 a_1250_231# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=3.024e+11p pd=2.4e+06u as=0p ps=0u
M1016 VGND a_341_93# a_299_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1880_119# a_1250_231# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_2037_442# a_2881_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1019 a_877_98# a_622_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1020 VPWR a_1250_231# a_1224_419# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1021 a_1250_231# a_1092_96# a_1418_125# VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=7.81e+11p ps=5.37e+06u
M1022 a_1418_125# a_1625_93# a_1250_231# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_2881_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1024 VPWR a_2037_442# a_1989_504# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 a_1418_125# SET_B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_2061_74# a_622_98# a_1881_420# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_2037_442# a_2881_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1028 a_221_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1029 a_1092_96# a_877_98# a_197_119# VPB pshort w=640000u l=180000u
+  ad=2.167e+11p pd=2.05e+06u as=3.52e+11p ps=3.66e+06u
M1030 a_1583_379# a_1092_96# a_1250_231# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1769_379# a_1250_231# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_341_93# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1033 a_197_119# SCE a_119_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1192_96# a_877_98# a_1092_96# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1035 a_2037_442# a_1881_420# a_2271_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1036 Q_N a_2037_442# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1037 a_1224_419# a_622_98# a_1092_96# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1092_96# a_622_98# a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_197_119# D a_221_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1989_504# a_877_98# a_1881_420# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_2387_392# a_1881_420# a_2037_442# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.7e+11p ps=2.74e+06u
M1042 a_27_464# a_341_93# a_197_119# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_341_93# SCE VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1044 VGND CLK a_622_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1045 a_2271_74# a_1625_93# a_2037_442# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_2037_442# SET_B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR RESET_B a_1625_93# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 Q a_2513_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=2.27097e+12p ps=1.957e+07u
M1001 VPWR SCD a_515_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.304e+11p ps=2e+06u
M1002 a_413_90# D a_312_90# VNB nlowvt w=420000u l=150000u
+  ad=3.26375e+11p pd=3.3e+06u as=1.491e+11p ps=1.55e+06u
M1003 VGND a_1747_74# a_2513_424# VNB nlowvt w=550000u l=150000u
+  ad=1.78918e+12p pd=1.476e+07u as=1.4575e+11p ps=1.63e+06u
M1004 a_1399_119# a_1369_93# a_1321_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1005 VGND a_2008_48# a_1966_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 VPWR a_1369_93# a_1331_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_1369_93# a_1235_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1008 VPWR a_1747_74# a_2513_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1009 a_2124_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 Q_N a_1747_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1011 a_413_90# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=4.654e+11p pd=5.04e+06u as=0p ps=0u
M1012 a_2008_48# a_1747_74# a_2124_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1013 VGND CLK a_819_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.54e+11p ps=2.22e+06u
M1014 a_1037_119# a_819_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1015 a_1747_74# a_819_119# a_1369_93# VPB pshort w=1e+06u l=180000u
+  ad=3.9355e+11p pd=3.45e+06u as=0p ps=0u
M1016 a_1966_74# a_819_119# a_1747_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.519e+11p ps=3.17e+06u
M1017 a_341_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1018 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=5.696e+11p ps=3.06e+06u
M1019 a_1235_119# a_1037_119# a_413_90# VPB pshort w=420000u l=180000u
+  ad=2.268e+11p pd=2.76e+06u as=0p ps=0u
M1020 a_2008_48# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1021 VPWR a_1747_74# a_2008_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_225_90# SCD a_545_97# VNB nlowvt w=420000u l=150000u
+  ad=2.64075e+11p pd=2.99e+06u as=8.82e+10p ps=1.26e+06u
M1023 a_312_90# a_27_74# a_225_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1331_463# a_819_119# a_1235_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR CLK a_819_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1026 Q_N a_1747_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1027 a_413_90# D a_341_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND RESET_B a_225_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1747_74# a_1037_119# a_1369_93# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1030 a_515_464# a_27_74# a_413_90# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1235_119# a_819_119# a_413_90# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1032 a_545_97# SCE a_413_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1972_489# a_1037_119# a_1747_74# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1034 VGND RESET_B a_1399_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1037_119# a_819_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1036 a_1321_119# a_1037_119# a_1235_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q a_2513_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1038 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1039 VPWR a_2008_48# a_1972_489# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1235_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1369_93# a_1235_119# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1370_290# a_1223_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=3.2444e+12p ps=2.643e+07u
M1001 VPWR a_2607_392# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1002 a_2000_74# a_852_119# a_1790_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.33e+11p ps=3.08e+06u
M1003 VGND RESET_B a_223_79# VNB nlowvt w=420000u l=150000u
+  ad=2.20072e+12p pd=1.854e+07u as=2.751e+11p ps=2.99e+06u
M1004 a_1790_74# a_852_119# a_1370_290# VPB pshort w=1e+06u l=180000u
+  ad=3.816e+11p pd=3.22e+06u as=0p ps=0u
M1005 Q_N a_1790_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 a_388_79# D a_310_464# VPB pshort w=640000u l=180000u
+  ad=6.96975e+11p pd=5.83e+06u as=1.536e+11p ps=1.76e+06u
M1007 a_1370_290# a_1223_119# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1008 VPWR a_1790_74# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR SCE a_27_79# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1010 a_2607_392# a_1790_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1011 VGND RESET_B a_1401_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1012 a_310_79# a_27_79# a_223_79# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1013 a_223_79# SCD a_547_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1014 a_1223_119# a_852_119# a_388_79# VNB nlowvt w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=3.906e+11p ps=3.54e+06u
M1015 a_1323_119# a_1025_119# a_1223_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1016 a_2006_373# a_1790_74# a_2158_74# VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1017 a_1790_74# a_1025_119# a_1370_290# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_2607_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1019 VPWR CLK a_852_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1020 VPWR a_1370_290# a_1328_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1021 VGND CLK a_852_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.95675e+11p ps=2.05e+06u
M1022 VPWR a_2006_373# a_1958_471# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1023 a_2006_373# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1024 a_2158_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q_N a_1790_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1026 a_388_79# D a_310_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_541_483# a_27_79# a_388_79# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1028 VPWR a_1790_74# a_2006_373# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_2607_392# a_1790_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1030 VGND SCE a_27_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1031 a_547_79# SCE a_388_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1223_119# a_1025_119# a_388_79# VPB pshort w=420000u l=180000u
+  ad=2.247e+11p pd=2.75e+06u as=0p ps=0u
M1033 a_1025_119# a_852_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1034 a_1223_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_388_79# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1025_119# a_852_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1037 VGND a_1790_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_2607_392# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_310_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1328_457# a_852_119# a_1223_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR SCD a_541_483# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1958_471# a_1025_119# a_1790_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1401_119# a_1370_290# a_1323_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 Q a_2607_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND a_2006_373# a_2000_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 VPWR CLK_N a_859_347# VPB pshort w=1e+06u l=180000u
+  ad=2.14562e+12p pd=1.792e+07u as=3.25e+11p ps=2.65e+06u
M1001 a_1273_131# a_859_347# a_287_464# VPB pshort w=420000u l=180000u
+  ad=2.268e+11p pd=2.76e+06u as=7.8e+11p ps=6.03e+06u
M1002 a_287_464# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND RESET_B a_1483_131# VNB nlowvt w=420000u l=150000u
+  ad=1.49337e+12p pd=1.266e+07u as=8.82e+10p ps=1.26e+06u
M1004 VGND a_2087_410# a_2073_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.05e+11p ps=1.34e+06u
M1005 a_2045_508# a_859_347# a_1827_144# VPB pshort w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=2.915e+11p ps=2.67e+06u
M1006 a_538_81# SCE a_287_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.465e+11p ps=3.33e+06u
M1007 VGND CLK_N a_859_347# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.442e+11p ps=2.14e+06u
M1008 a_1069_74# a_859_347# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.257e+11p pd=2.09e+06u as=0p ps=0u
M1009 a_2265_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1010 a_2087_410# a_1827_144# a_2265_74# VNB nlowvt w=420000u l=150000u
+  ad=2.1e+11p pd=1.84e+06u as=0p ps=0u
M1011 VPWR SCE a_27_88# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1012 a_209_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1013 VPWR a_2087_410# a_2045_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q a_2492_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1015 a_474_464# a_27_88# a_287_464# VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1016 a_1483_131# a_1417_294# a_1409_131# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=9.24e+10p ps=1.28e+06u
M1017 Q a_2492_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1018 a_324_81# a_27_88# a_239_81# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1019 a_2087_410# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1020 a_287_464# D a_324_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1273_131# a_1069_74# a_287_464# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1022 VPWR a_1827_144# a_2087_410# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND RESET_B a_239_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1381_457# a_1069_74# a_1273_131# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1025 VPWR a_1827_144# a_2492_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1026 a_2073_74# a_1069_74# a_1827_144# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=6.59025e+11p ps=4.26e+06u
M1027 VGND a_1827_144# a_2492_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1028 a_1409_131# a_859_347# a_1273_131# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1069_74# a_859_347# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1030 a_1273_131# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1827_144# a_1069_74# a_1417_294# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.55e+11p ps=3.51e+06u
M1032 a_239_81# SCD a_538_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1417_294# a_1381_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_287_464# D a_209_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1417_294# a_1273_131# VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=2.4e+06u as=0p ps=0u
M1036 VPWR SCD a_474_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND SCE a_27_88# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1038 a_1417_294# a_1273_131# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1827_144# a_859_347# a_1417_294# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1234_119# a_1037_387# a_303_464# VPB pshort w=420000u l=180000u
+  ad=2.576e+11p pd=2.93e+06u as=9.24e+11p ps=6.48e+06u
M1001 a_1320_119# a_1037_387# a_1234_119# VNB nlowvt w=420000u l=150000u
+  ad=9.87e+10p pd=1.31e+06u as=1.176e+11p ps=1.4e+06u
M1002 a_219_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=2.08418e+12p ps=1.846e+07u
M1003 VGND a_1997_272# a_1972_74# VNB nlowvt w=420000u l=150000u
+  ad=1.60052e+12p pd=1.375e+07u as=8.82e+10p ps=1.26e+06u
M1004 a_1972_74# a_835_93# a_1745_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.687e+11p ps=3.25e+06u
M1005 VPWR SCE a_27_88# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 a_1745_74# a_1037_387# a_1367_93# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1007 Q a_2402_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 a_312_81# a_27_88# a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.499e+11p ps=2.87e+06u
M1009 a_303_464# D a_312_81# VNB nlowvt w=420000u l=150000u
+  ad=3.738e+11p pd=3.46e+06u as=0p ps=0u
M1010 a_1234_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_2402_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1012 VGND RESET_B a_1397_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_303_464# D a_219_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1996_508# a_1037_387# a_1745_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=4.21675e+11p ps=3.58e+06u
M1015 a_225_81# SCD a_545_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 a_535_464# a_27_88# a_303_464# VPB pshort w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1017 a_1346_461# a_835_93# a_1234_119# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 VPWR CLK a_835_93# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1019 VPWR SCD a_535_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1397_119# a_1367_93# a_1320_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1997_272# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1022 a_1997_272# a_1745_74# a_2135_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1023 a_303_464# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1745_74# a_1997_272# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_545_81# SCE a_303_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1367_93# a_1234_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1027 a_2402_424# a_1745_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1028 VPWR a_1367_93# a_1346_461# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND CLK a_835_93# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.8265e+11p ps=2.43e+06u
M1030 a_1037_387# a_835_93# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1031 a_1745_74# a_835_93# a_1367_93# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1037_387# a_835_93# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1033 a_1367_93# a_1234_119# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SCE a_27_88# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1035 a_1234_119# a_835_93# a_303_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND RESET_B a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_1997_272# a_1996_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_2135_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2402_424# a_1745_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_390_81# D a_343_483# VPB pshort w=640000u l=180000u
+  ad=5.4e+11p pd=5.28e+06u as=1.472e+11p ps=1.74e+06u
M1001 VPWR a_2495_392# Q VPB pshort w=1.12e+06u l=180000u
+  ad=2.9811e+12p pd=2.35e+07u as=3.024e+11p ps=2.78e+06u
M1002 a_1235_119# a_1037_119# a_390_81# VPB pshort w=420000u l=180000u
+  ad=2.394e+11p pd=2.82e+06u as=0p ps=0u
M1003 Q a_2495_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.0718e+12p ps=1.661e+07u
M1004 VGND RESET_B a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.88e+06u
M1005 VPWR a_2082_446# a_2040_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_1383_349# a_1235_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=4.6755e+11p pd=3.07e+06u as=0p ps=0u
M1007 VGND RESET_B a_1432_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 a_547_81# SCE a_390_81# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.927e+11p ps=3.55e+06u
M1009 a_2078_74# a_837_119# a_1824_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=5.504e+11p ps=3.72e+06u
M1010 VGND a_2082_446# a_2078_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1012 a_343_483# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1235_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_312_81# a_27_74# a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1015 a_390_81# D a_312_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND CLK a_837_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.0225e+11p ps=2.04e+06u
M1017 a_1037_119# a_837_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1018 a_2082_446# a_1824_74# a_2242_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1019 a_2082_446# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1020 a_1824_74# a_837_119# a_1383_349# VPB pshort w=1e+06u l=180000u
+  ad=4.2595e+11p pd=3.6e+06u as=0p ps=0u
M1021 a_2040_508# a_1037_119# a_1824_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1432_119# a_1383_349# a_1354_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1023 a_390_81# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1824_74# a_2082_446# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1339_457# a_837_119# a_1235_119# VPB pshort w=420000u l=180000u
+  ad=9.24e+10p pd=1.28e+06u as=0p ps=0u
M1026 a_2242_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR CLK a_837_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1028 a_1824_74# a_1037_119# a_1383_349# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.627e+11p ps=2.19e+06u
M1029 a_2495_392# a_1824_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1030 VGND a_2495_392# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1235_119# a_837_119# a_390_81# VNB nlowvt w=420000u l=150000u
+  ad=1.869e+11p pd=1.73e+06u as=0p ps=0u
M1032 a_1354_119# a_1037_119# a_1235_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1383_349# a_1339_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1037_119# a_837_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1035 a_225_81# SCD a_547_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_2495_392# a_1824_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1038 a_517_483# a_27_74# a_390_81# VPB pshort w=640000u l=180000u
+  ad=2.304e+11p pd=2e+06u as=0p ps=0u
M1039 VPWR SCD a_517_483# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1383_349# a_1235_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Q a_2495_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1397_138# a_1367_112# a_1319_138# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1001 VPWR a_1745_74# a_2339_74# VPB pshort w=840000u l=180000u
+  ad=3.24455e+12p pd=2.618e+07u as=2.268e+11p ps=2.22e+06u
M1002 VPWR a_1367_112# a_1345_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1003 a_1233_138# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=2.52e+11p pd=2.88e+06u as=0p ps=0u
M1004 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1005 a_225_81# SCD a_555_81# VNB nlowvt w=420000u l=150000u
+  ad=2.583e+11p pd=2.91e+06u as=8.82e+10p ps=1.26e+06u
M1006 a_1745_74# a_1037_387# a_1367_112# VNB nlowvt w=640000u l=150000u
+  ad=4.33e+11p pd=3.08e+06u as=2.33e+11p ps=2.13e+06u
M1007 a_312_81# a_27_74# a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
M1008 a_415_81# D a_312_81# VNB nlowvt w=420000u l=150000u
+  ad=3.423e+11p pd=3.31e+06u as=0p ps=0u
M1009 VGND a_2339_74# Q VNB nlowvt w=740000u l=150000u
+  ad=2.376e+12p pd=1.764e+07u as=4.144e+11p ps=4.08e+06u
M1010 VPWR a_2003_48# a_1985_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1011 VGND a_1745_74# a_2339_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1012 a_1345_463# a_834_93# a_1233_138# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND RESET_B a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1985_508# a_1037_387# a_1745_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=4.06975e+11p ps=3.51e+06u
M1015 Q a_2339_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1016 a_1233_138# a_1037_387# a_415_81# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=4.728e+11p ps=5.07e+06u
M1017 a_1319_138# a_1037_387# a_1233_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1018 a_1367_112# a_1233_138# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1019 VPWR a_2339_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q a_2339_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_415_81# D a_343_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1022 a_1745_74# a_834_93# a_1367_112# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_2339_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_517_464# a_27_74# a_415_81# VPB pshort w=640000u l=180000u
+  ad=2.432e+11p pd=2.04e+06u as=0p ps=0u
M1025 a_555_81# SCE a_415_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR CLK a_834_93# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1027 a_1233_138# a_834_93# a_415_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1367_112# a_1233_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2339_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_2003_48# a_1745_74# a_2141_74# VNB nlowvt w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=8.82e+10p ps=1.26e+06u
M1031 a_2003_48# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.491e+11p pd=1.55e+06u as=0p ps=0u
M1032 VGND a_2003_48# a_1955_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1033 Q a_2339_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND RESET_B a_1397_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_415_81# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1955_74# a_834_93# a_1745_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_2339_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND CLK a_834_93# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.7955e+11p ps=2.44e+06u
M1039 a_343_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1037_387# a_834_93# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1041 a_1037_387# a_834_93# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.924e+11p pd=2e+06u as=0p ps=0u
M1042 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1043 VPWR SCD a_517_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR a_1745_74# a_2003_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_2141_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_2339_74# a_1745_74# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 Q_N a_1762_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=1.9498e+12p ps=1.823e+07u
M1001 a_1411_74# a_995_74# a_1163_48# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1002 a_419_464# a_27_74# a_293_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=4.014e+11p ps=3.56e+06u
M1003 a_1876_74# a_594_74# a_1762_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.391e+11p ps=2.12e+06u
M1004 a_1954_74# a_1924_48# a_1876_74# VNB nlowvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1005 VGND a_1163_48# a_1115_74# VNB nlowvt w=420000u l=150000u
+  ad=2.17215e+12p pd=1.688e+07u as=1.008e+11p ps=1.32e+06u
M1006 a_1924_48# a_1762_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1007 a_1115_74# a_781_74# a_995_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.89e+11p ps=1.74e+06u
M1008 a_1603_347# a_594_74# a_1762_74# VPB pshort w=1e+06u l=180000u
+  ad=5.5e+11p pd=5.1e+06u as=4.117e+11p ps=4.11e+06u
M1009 Q_N a_1762_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1011 a_209_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1012 VGND SET_B a_1954_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR SCD a_419_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND SET_B a_1411_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_392_74# SCE a_293_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.0425e+11p ps=3.2e+06u
M1016 VGND SCD a_392_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_293_464# D a_209_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1762_74# a_2556_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1019 a_781_74# a_594_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1020 a_1136_478# a_594_74# a_995_74# VPB pshort w=420000u l=180000u
+  ad=1.548e+11p pd=1.67e+06u as=1.99125e+11p ps=1.84e+06u
M1021 VPWR a_1163_48# a_1136_478# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_995_74# a_781_74# a_293_464# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK a_594_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1024 a_1684_74# a_995_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1025 a_1762_74# a_781_74# a_1684_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR CLK a_594_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1027 Q a_2556_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1028 VPWR a_1924_48# a_1712_374# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.618e+11p ps=4.39e+06u
M1029 VPWR a_1762_74# a_1924_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1030 a_781_74# a_594_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1031 Q a_2556_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1032 a_1762_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1762_74# a_781_74# a_1712_374# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_1762_74# a_2556_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1035 VPWR SET_B a_1163_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.722e+11p ps=1.66e+06u
M1036 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_995_74# a_594_74# a_293_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1163_48# a_995_74# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_228_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1040 a_293_464# D a_228_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1603_347# a_995_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_2067_74# a_3177_368# VPB pshort w=1e+06u l=180000u
+  ad=3.4604e+12p pd=2.71e+07u as=2.8e+11p ps=2.56e+06u
M1001 VGND a_3177_368# Q VNB nlowvt w=740000u l=150000u
+  ad=2.2419e+12p pd=2.069e+07u as=2.072e+11p ps=2.04e+06u
M1002 a_1204_463# a_619_368# a_1069_81# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.344e+11p ps=1.48e+06u
M1003 a_1789_424# a_1069_81# VPWR VPB pshort w=840000u l=180000u
+  ad=7.392e+11p pd=6.8e+06u as=0p ps=0u
M1004 Q_N a_2067_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VGND a_1069_81# a_1794_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=6.208e+11p ps=5.78e+06u
M1006 a_1069_81# a_871_74# a_307_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.672e+11p ps=3.46e+06u
M1007 a_223_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1008 a_2501_74# a_619_368# a_2067_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=5.999e+11p ps=4.61e+06u
M1009 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1010 a_2067_74# a_871_74# a_2277_455# VPB pshort w=420000u l=180000u
+  ad=4.62e+11p pd=5.02e+06u as=2.373e+11p ps=2.81e+06u
M1011 a_1794_74# a_1069_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_2067_74# a_3177_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1013 a_1567_74# a_1069_81# a_1252_376# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1014 VGND SET_B a_1567_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND SCD a_495_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 VPWR a_2513_258# a_2277_455# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_495_74# SCE a_307_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.515e+11p ps=3.83e+06u
M1018 a_2067_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1069_81# a_619_368# a_307_74# VNB nlowvt w=420000u l=150000u
+  ad=3.675e+11p pd=2.59e+06u as=0p ps=0u
M1020 a_2579_74# a_2513_258# a_2501_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1021 VGND SET_B a_2579_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q a_3177_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_2067_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.22e+11p pd=2.08e+06u as=0p ps=0u
M1024 VGND a_1252_376# a_1274_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VGND a_2067_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1274_81# a_871_74# a_1069_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_421_464# a_27_74# a_307_74# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1028 a_2067_74# a_619_368# a_1789_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2067_74# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1252_376# a_1204_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1789_424# a_619_368# a_2067_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1794_74# a_871_74# a_2067_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_307_74# D a_223_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR SET_B a_1252_376# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.554e+11p ps=1.58e+06u
M1035 a_871_74# a_619_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1036 VPWR CLK a_619_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1037 a_229_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1038 a_307_74# D a_229_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2067_74# a_871_74# a_1794_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_2513_258# a_2067_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1041 VPWR SCD a_421_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1252_376# a_1069_81# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND CLK a_619_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1044 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1045 VPWR a_2067_74# a_2513_258# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1046 a_871_74# a_619_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.528e+11p pd=2.87e+06u as=0p ps=0u
M1047 Q a_3177_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1048 VPWR a_1069_81# a_1789_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR a_3177_368# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 a_1686_74# a_998_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.66425e+12p ps=1.358e+07u
M1001 a_1764_74# a_800_74# a_1686_74# VNB nlowvt w=640000u l=150000u
+  ad=3.547e+11p pd=2.44e+06u as=0p ps=0u
M1002 a_998_81# a_800_74# a_292_464# VPB pshort w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=4.056e+11p ps=3.58e+06u
M1003 a_238_74# a_27_464# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1004 VGND SCD a_402_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 a_402_74# SCE a_292_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.373e+11p ps=2.81e+06u
M1006 VGND CLK a_599_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1007 a_1613_341# a_998_81# VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.35e+11p pd=5.07e+06u as=2.003e+12p ps=1.815e+07u
M1008 a_1988_74# a_1958_48# a_1910_74# VNB nlowvt w=420000u l=150000u
+  ad=3.192e+11p pd=2.36e+06u as=1.008e+11p ps=1.32e+06u
M1009 VGND a_1198_55# a_1150_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 a_1131_457# a_599_74# a_998_81# VPB pshort w=420000u l=180000u
+  ad=1.407e+11p pd=1.51e+06u as=0p ps=0u
M1011 a_1150_81# a_800_74# a_998_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.562e+11p ps=2.06e+06u
M1012 VGND SET_B a_1426_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_418_464# a_27_464# a_292_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1014 a_998_81# a_599_74# a_292_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_800_74# a_599_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 a_1613_341# a_599_74# a_1764_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.18e+11p ps=4.14e+06u
M1017 VPWR SCE a_27_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1018 a_208_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 VPWR SCD a_418_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1198_55# a_1131_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q a_2395_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1022 VGND SET_B a_1988_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_2395_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1024 VPWR SET_B a_1198_55# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1025 VGND SCE a_27_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1026 VPWR a_1958_48# a_1721_374# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.655e+11p ps=4.42e+06u
M1027 VPWR a_1764_74# a_2395_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1028 a_292_464# D a_208_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR CLK a_599_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1030 a_1198_55# a_998_81# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1764_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1426_118# a_998_81# a_1198_55# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 a_800_74# a_599_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.908e+11p pd=2.8e+06u as=0p ps=0u
M1034 a_292_464# D a_238_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_1764_74# a_1958_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1036 VGND a_1764_74# a_2395_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=3.85e+11p ps=2.5e+06u
M1037 a_1910_74# a_599_74# a_1764_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1764_74# a_800_74# a_1721_374# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1958_48# a_1764_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 a_1587_379# a_991_81# VPWR VPB pshort w=840000u l=180000u
+  ad=4.536e+11p pd=4.44e+06u as=2.366e+12p ps=2.199e+07u
M1001 a_1804_424# a_795_74# a_1641_74# VNB nlowvt w=640000u l=150000u
+  ad=4.292e+11p pd=3.97e+06u as=3.584e+11p ps=3.68e+06u
M1002 VPWR a_1804_424# a_2611_98# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1003 a_1587_379# a_608_74# a_1804_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=7.287e+11p ps=6.51e+06u
M1004 VPWR a_2611_98# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1005 a_419_464# a_27_74# a_293_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=4.056e+11p ps=3.58e+06u
M1006 a_795_74# a_608_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.0955e+12p ps=1.834e+07u
M1007 VPWR a_991_81# a_1587_379# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_2186_367# a_2144_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 VPWR a_1804_424# a_2186_367# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1010 a_1804_424# a_608_74# a_1587_379# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1185_55# a_991_81# VPWR VPB pshort w=420000u l=180000u
+  ad=1.323e+11p pd=1.47e+06u as=0p ps=0u
M1012 VGND CLK a_608_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1013 a_1804_424# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q a_2611_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1015 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1016 a_209_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1017 VPWR SCD a_419_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1120_483# a_608_74# a_991_81# VPB pshort w=420000u l=180000u
+  ad=1.588e+11p pd=1.72e+06u as=1.7185e+11p ps=1.81e+06u
M1019 a_2144_508# a_795_74# a_1804_424# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1185_55# a_1143_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1021 VPWR SET_B a_1185_55# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1804_424# a_2611_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1023 a_293_464# D a_209_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_991_81# a_608_74# a_293_464# VNB nlowvt w=420000u l=150000u
+  ad=2.562e+11p pd=2.06e+06u as=2.352e+11p ps=2.8e+06u
M1025 VGND SET_B a_2219_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1026 a_1429_74# a_991_81# a_1185_55# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1027 VGND SET_B a_1429_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_293_464# D a_239_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1029 a_1641_74# a_991_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_2186_367# a_1804_424# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1031 a_1143_81# a_795_74# a_991_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR CLK a_608_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1033 VGND a_991_81# a_1641_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_991_81# a_795_74# a_293_464# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND SCD a_403_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1036 a_1641_74# a_795_74# a_1804_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_2611_98# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_239_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_403_74# SCE a_293_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_795_74# a_608_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.908e+11p pd=2.8e+06u as=0p ps=0u
M1041 a_2219_74# a_2186_367# a_2141_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1042 VPWR a_1185_55# a_1120_483# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1044 a_2141_74# a_608_74# a_1804_424# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 Q a_2611_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 Q a_2580_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=2.9103e+12p ps=2.649e+07u
M1001 Q a_2580_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=5.291e+11p pd=4.39e+06u as=2.27325e+12p ps=1.996e+07u
M1002 a_1017_81# a_616_74# a_291_464# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=3.592e+11p ps=3.44e+06u
M1003 VGND SET_B a_1445_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 a_2227_74# a_2191_180# a_2149_74# VNB nlowvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.008e+11p ps=1.32e+06u
M1005 VGND a_1823_524# a_2580_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1006 a_1823_524# a_803_74# a_1677_74# VNB nlowvt w=640000u l=150000u
+  ad=3.963e+11p pd=3.85e+06u as=3.584e+11p ps=3.68e+06u
M1007 VPWR a_2191_180# a_2106_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.869e+11p ps=1.73e+06u
M1008 a_1017_81# a_803_74# a_291_464# VPB pshort w=420000u l=180000u
+  ad=1.8235e+11p pd=1.93e+06u as=4.056e+11p ps=3.58e+06u
M1009 a_2580_74# a_1823_524# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1010 VPWR a_1201_55# a_1143_495# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.6975e+11p ps=1.87e+06u
M1011 a_1823_524# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=5.793e+11p pd=5.97e+06u as=0p ps=0u
M1012 VGND a_1017_81# a_1677_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1143_495# a_616_74# a_1017_81# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_1823_524# a_2580_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_2580_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_417_74# SCE a_291_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1017 VGND SCD a_417_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1201_55# a_1153_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 a_1153_81# a_803_74# a_1017_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_803_74# a_616_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 VGND a_2580_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1445_74# a_1017_81# a_1201_55# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1023 VPWR SET_B a_1201_55# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1024 a_1623_373# a_1017_81# VPWR VPB pshort w=840000u l=180000u
+  ad=4.536e+11p pd=4.44e+06u as=0p ps=0u
M1025 VGND CLK a_616_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 a_2149_74# a_616_74# a_1823_524# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_417_464# a_27_74# a_291_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1028 a_1201_55# a_1017_81# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1017_81# a_1623_373# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_2580_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_2580_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2106_508# a_803_74# a_1823_524# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1034 a_207_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1035 VPWR SCD a_417_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1677_74# a_803_74# a_1823_524# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_1823_524# a_2191_180# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1038 VGND SET_B a_2227_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2191_180# a_1823_524# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1040 a_222_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1041 a_291_464# D a_222_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR CLK a_616_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1043 a_1623_373# a_616_74# a_1823_524# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_291_464# D a_207_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1046 Q a_2580_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_1823_524# a_616_74# a_1623_373# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_803_74# a_616_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.088e+11p pd=2.9e+06u as=0p ps=0u
M1049 a_1677_74# a_1017_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VPWR a_2580_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1529_74# a_612_74# a_1243_398# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=6.216e+11p ps=3.16e+06u
M1001 a_1723_48# a_1529_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=1.8401e+12p ps=1.538e+07u
M1002 VPWR a_1723_48# a_1694_508# VPB pshort w=420000u l=180000u
+  ad=2.5456e+12p pd=2.012e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_434_74# SCE a_296_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.423e+11p ps=3.31e+06u
M1004 VPWR a_1723_48# a_2216_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1005 Q a_1723_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1006 a_1157_100# a_828_74# a_1021_100# VNB nlowvt w=420000u l=150000u
+  ad=1.932e+11p pd=1.76e+06u as=2.226e+11p ps=1.9e+06u
M1007 a_218_74# a_31_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1008 a_296_74# D a_218_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR SCD a_410_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.304e+11p ps=2e+06u
M1010 a_1529_74# a_828_74# a_1243_398# VNB nlowvt w=550000u l=150000u
+  ad=2.887e+11p pd=2.32e+06u as=1.5675e+11p ps=1.67e+06u
M1011 a_1243_398# a_1021_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q a_1723_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 a_612_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1014 a_1723_48# a_1529_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1015 a_828_74# a_612_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1016 VGND a_1243_398# a_1157_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1681_74# a_612_74# a_1529_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1018 a_236_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_1243_398# a_1021_100# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1694_508# a_828_74# a_1529_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1723_48# a_1681_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR SCE a_31_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1023 a_612_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1024 VGND SCE a_31_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1025 a_828_74# a_612_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1026 Q_N a_2216_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1027 VGND SCD a_434_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_296_74# D a_236_464# VPB pshort w=640000u l=180000u
+  ad=2.841e+11p pd=3.19e+06u as=0p ps=0u
M1029 a_1021_100# a_828_74# a_296_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1030 a_1021_100# a_612_74# a_296_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_1243_398# a_1183_496# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1032 a_410_464# a_31_74# a_296_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1183_496# a_612_74# a_1021_100# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q_N a_2216_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1035 VGND a_1723_48# a_2216_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 VGND a_1711_48# Q VNB nlowvt w=740000u l=150000u
+  ad=2.2043e+12p pd=1.954e+07u as=2.072e+11p ps=2.04e+06u
M1001 a_1511_74# a_630_74# a_1243_48# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=5.166e+11p ps=2.91e+06u
M1002 VGND a_2322_368# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.183e+11p ps=2.07e+06u
M1003 VPWR a_1711_48# a_1694_508# VPB pshort w=420000u l=180000u
+  ad=3.0047e+12p pd=2.544e+07u as=1.008e+11p ps=1.32e+06u
M1004 VPWR SCE a_36_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.336e+11p ps=2.01e+06u
M1005 a_630_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 a_241_453# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1007 a_630_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=5.488e+11p pd=3.22e+06u as=0p ps=0u
M1008 a_1220_499# a_630_74# a_1021_97# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.491e+11p ps=1.55e+06u
M1009 Q a_1711_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1010 VPWR a_1711_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_1243_48# a_1220_499# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1663_74# a_630_74# a_1511_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.887e+11p ps=2.32e+06u
M1013 VGND a_1711_48# a_1663_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1711_48# a_1511_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1015 a_828_74# a_630_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1016 a_301_74# D a_241_453# VPB pshort w=640000u l=180000u
+  ad=3.256e+11p pd=3.33e+06u as=0p ps=0u
M1017 a_223_74# a_36_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_301_74# D a_223_74# VNB nlowvt w=420000u l=150000u
+  ad=3.654e+11p pd=3.42e+06u as=0p ps=0u
M1019 a_1243_48# a_1021_97# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1243_48# a_1173_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.6425e+11p ps=1.77e+06u
M1021 a_426_453# a_36_74# a_301_74# VPB pshort w=640000u l=180000u
+  ad=1.952e+11p pd=1.89e+06u as=0p ps=0u
M1022 a_1694_508# a_828_74# a_1511_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1021_97# a_828_74# a_301_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1021_97# a_630_74# a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=2.562e+11p pd=2.06e+06u as=0p ps=0u
M1025 a_1243_48# a_1021_97# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=0p ps=0u
M1026 Q_N a_2322_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1711_48# a_2322_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1028 a_828_74# a_630_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1029 Q a_1711_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1711_48# a_2322_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1031 VGND SCD a_450_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1032 a_1711_48# a_1511_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1033 a_450_74# SCE a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q_N a_2322_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1035 a_1173_97# a_828_74# a_1021_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_2322_368# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR SCD a_426_453# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND SCE a_36_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1039 a_1511_74# a_828_74# a_1243_48# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_1520_74# a_828_74# a_1239_74# VNB nlowvt w=550000u l=150000u
+  ad=3.223e+11p pd=2.48e+06u as=1.5675e+11p ps=1.67e+06u
M1001 Q a_1736_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=2.1858e+12p ps=1.697e+07u
M1002 VPWR SCD a_415_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.304e+11p ps=2e+06u
M1003 a_630_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.52935e+12p ps=1.307e+07u
M1004 a_630_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 VGND a_1736_74# a_1688_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VGND SCE a_35_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1007 a_1018_100# a_630_74# a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=3.612e+11p ps=3.4e+06u
M1008 a_828_74# a_630_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1009 a_1736_74# a_1520_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.4575e+11p pd=1.63e+06u as=0p ps=0u
M1010 a_1691_508# a_828_74# a_1520_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=3.738e+11p ps=2.73e+06u
M1011 a_1239_74# a_1018_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_241_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1013 a_1205_508# a_630_74# a_1018_100# VPB pshort w=420000u l=180000u
+  ad=9.24e+10p pd=1.28e+06u as=1.344e+11p ps=1.48e+06u
M1014 VPWR SCE a_35_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1015 a_1018_100# a_828_74# a_301_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.904e+11p ps=3.22e+06u
M1016 a_1239_74# a_1018_100# VPWR VPB pshort w=840000u l=180000u
+  ad=4.41e+11p pd=2.73e+06u as=0p ps=0u
M1017 Q a_1736_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=0p ps=0u
M1018 a_828_74# a_630_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1019 VPWR a_1239_74# a_1205_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_223_74# a_35_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1021 a_301_74# D a_223_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1736_74# a_1691_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1688_100# a_630_74# a_1520_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_1239_74# a_1154_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.785e+11p ps=1.69e+06u
M1025 a_301_74# D a_241_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1520_74# a_630_74# a_1239_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_415_464# a_35_74# a_301_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND SCD a_450_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1029 a_450_74# SCE a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1154_100# a_828_74# a_1018_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1736_74# a_1520_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_1707_496# a_846_74# a_1595_424# VPB pshort w=420000u l=180000u
+  ad=2.562e+11p pd=2.06e+06u as=2.754e+11p ps=2.44e+06u
M1001 a_1044_100# a_634_74# a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=3.045e+11p pd=2.29e+06u as=3.528e+11p ps=3.36e+06u
M1002 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=2.72693e+12p pd=2.061e+07u as=1.792e+11p ps=1.84e+06u
M1003 a_1595_424# a_634_74# a_1287_320# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.2e+11p ps=2.68e+06u
M1004 VGND SCD a_442_74# VNB nlowvt w=420000u l=150000u
+  ad=1.84785e+12p pd=1.542e+07u as=1.008e+11p ps=1.32e+06u
M1005 VGND a_1829_398# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.13e+06u
M1006 a_301_74# D a_219_453# VPB pshort w=640000u l=180000u
+  ad=4.472e+11p pd=3.71e+06u as=1.536e+11p ps=1.76e+06u
M1007 a_1219_100# a_846_74# a_1044_100# VNB nlowvt w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=0p ps=0u
M1008 a_1287_320# a_1044_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=3.795e+11p pd=2.48e+06u as=0p ps=0u
M1009 a_1829_398# a_1595_424# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1010 VGND a_1287_320# a_1219_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1595_424# a_846_74# a_1287_320# VNB nlowvt w=550000u l=150000u
+  ad=1.8825e+11p pd=1.82e+06u as=0p ps=0u
M1012 a_634_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1013 a_442_74# SCE a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_1829_398# a_1707_496# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_223_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1016 a_301_74# D a_223_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1829_398# a_1595_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1018 VPWR SCD a_442_453# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1019 a_846_74# a_634_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1020 VPWR a_1287_320# a_1213_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.554e+11p ps=1.58e+06u
M1021 a_1787_74# a_634_74# a_1595_424# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1022 VGND a_1829_398# a_1787_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1044_100# a_846_74# a_301_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1024 Q a_1829_398# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1213_508# a_634_74# a_1044_100# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_1829_398# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 a_1287_320# a_1044_100# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_1829_398# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_442_453# a_27_74# a_301_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_846_74# a_634_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1031 a_634_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1032 a_219_453# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 VPWR SCD a_415_464# VPB pshort w=640000u l=180000u
+  ad=2.83978e+12p pd=2.238e+07u as=2.304e+11p ps=2e+06u
M1001 a_630_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_1026_100# a_828_74# a_301_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=2.904e+11p ps=3.22e+06u
M1003 a_630_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.77695e+12p ps=1.604e+07u
M1004 VGND a_1814_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.773e+11p ps=4.25e+06u
M1005 Q a_1814_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1006 a_1217_506# a_630_74# a_1026_100# VPB pshort w=420000u l=180000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1007 VPWR a_1814_48# a_1767_476# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VPWR a_1587_74# a_1814_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1009 VPWR a_1257_74# a_1217_506# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND SCD a_452_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1011 a_452_74# SCE a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.738e+11p ps=3.46e+06u
M1012 a_1162_100# a_828_74# a_1026_100# VNB nlowvt w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=2.226e+11p ps=1.9e+06u
M1013 a_241_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1014 VPWR a_1814_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR SCE a_36_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1016 Q a_1814_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q a_1814_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1814_48# a_1766_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 Q a_1814_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1766_74# a_630_74# a_1587_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4e+11p ps=2.59e+06u
M1021 a_828_74# a_630_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_223_74# a_36_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1023 a_301_74# D a_223_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1814_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_828_74# a_630_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1026 a_301_74# D a_241_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1026_100# a_630_74# a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1814_48# a_1587_74# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_415_464# a_36_74# a_301_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_1587_74# a_1814_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1031 VGND a_1814_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1587_74# a_828_74# a_1257_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.365e+11p ps=1.96e+06u
M1033 a_1587_74# a_630_74# a_1257_74# VPB pshort w=840000u l=180000u
+  ad=2.709e+11p pd=2.4e+06u as=7.308e+11p ps=3.42e+06u
M1034 VGND a_1257_74# a_1162_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1257_74# a_1026_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCE a_36_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_1257_74# a_1026_100# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1767_476# a_828_74# a_1587_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_114_112# GATE a_119_424# VPB pshort w=840000u l=180000u
+  ad=4.704e+11p pd=4.48e+06u as=1.764e+11p ps=2.1e+06u
M1001 a_709_54# a_566_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.81885e+12p ps=1.43e+07u
M1002 a_725_492# a_288_48# a_566_74# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=2.92075e+11p ps=2.68e+06u
M1003 a_318_74# a_288_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.3368e+12p ps=1.136e+07u
M1004 a_1238_94# CLK VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1005 VGND CLK a_288_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1006 a_1166_94# CLK VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1007 a_1238_94# a_709_54# a_1166_94# VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1008 a_119_424# SCE VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_709_54# a_1238_94# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_709_54# a_566_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1011 a_566_74# a_318_74# a_114_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND GATE a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=4.4825e+11p ps=3.83e+06u
M1013 a_114_112# SCE VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 GCLK a_1238_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=4.088e+11p pd=2.97e+06u as=0p ps=0u
M1015 a_667_80# a_318_74# a_566_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.846e+11p ps=1.81e+06u
M1016 VGND a_709_54# a_667_80# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_566_74# a_288_48# a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_709_54# a_725_492# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 GCLK a_1238_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1020 VPWR CLK a_288_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1021 a_318_74# a_288_48# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_706_317# a_580_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=2.04535e+12p ps=1.691e+07u
M1001 GCLK a_1198_374# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1002 VGND CLK a_288_48# VNB nlowvt w=740000u l=150000u
+  ad=1.5071e+12p pd=1.328e+07u as=2.109e+11p ps=2.05e+06u
M1003 VPWR a_1198_374# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_706_317# a_580_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_580_74# a_318_74# a_114_112# VPB pshort w=840000u l=180000u
+  ad=2.583e+11p pd=2.37e+06u as=4.536e+11p ps=4.44e+06u
M1006 a_318_74# a_288_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VPWR a_706_317# a_711_451# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1008 a_114_112# GATE a_117_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1009 GCLK a_1198_374# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1010 VPWR CLK a_288_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1011 a_1198_374# a_706_317# a_1198_74# VNB nlowvt w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=1.554e+11p ps=1.9e+06u
M1012 a_318_74# a_288_48# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1013 a_711_451# a_288_48# a_580_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND GATE a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=4.8675e+11p ps=3.97e+06u
M1015 a_114_112# SCE VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1198_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_1198_374# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_685_81# a_318_74# a_580_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.9475e+11p ps=1.85e+06u
M1019 VGND a_706_317# a_685_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_706_317# a_1198_374# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.85e+11p ps=2.97e+06u
M1021 a_1198_374# CLK VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_424# SCE VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_580_74# a_288_48# a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 VGND a_1292_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=1.98545e+12p pd=1.63e+07u as=4.514e+11p ps=4.18e+06u
M1001 a_119_143# GATE a_119_395# VPB pshort w=840000u l=180000u
+  ad=4.704e+11p pd=4.48e+06u as=2.016e+11p ps=2.16e+06u
M1002 VPWR CLK a_324_79# VPB pshort w=840000u l=180000u
+  ad=2.4738e+12p pd=1.955e+07u as=2.394e+11p ps=2.25e+06u
M1003 VGND a_1292_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_354_105# a_324_79# VPWR VPB pshort w=840000u l=180000u
+  ad=3.907e+11p pd=2.99e+06u as=0p ps=0u
M1005 a_634_74# a_354_105# a_119_143# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=0p ps=0u
M1006 a_792_48# a_634_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VGND a_792_48# a_744_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 a_788_455# a_324_79# a_634_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 GCLK a_1292_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=8.008e+11p pd=5.91e+06u as=0p ps=0u
M1010 VPWR a_1292_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1292_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1012 a_1292_368# a_792_48# a_1292_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 VGND CLK a_324_79# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1014 VPWR a_792_48# a_788_455# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 GCLK a_1292_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_1292_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_744_74# a_354_105# a_634_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.1025e+11p ps=1.9e+06u
M1018 GCLK a_1292_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_792_48# a_1292_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.208e+11p ps=3.17e+06u
M1020 a_1292_368# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_354_105# a_324_79# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_792_48# a_634_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1023 a_119_143# SCE VGND VNB nlowvt w=550000u l=150000u
+  ad=5.61e+11p pd=4.24e+06u as=0p ps=0u
M1024 a_634_74# a_324_79# a_119_143# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_119_395# SCE VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND GATE a_119_143# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 GCLK a_1292_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1549_74# a_1351_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=2.80005e+12p ps=2.337e+07u
M1001 a_1747_118# a_1351_74# a_697_113# VNB nlowvt w=420000u l=150000u
+  ad=2.478e+11p pd=2.02e+06u as=3.885e+11p ps=4.37e+06u
M1002 a_1895_118# a_1549_74# a_1747_118# VNB nlowvt w=420000u l=150000u
+  ad=1.617e+11p pd=1.61e+06u as=0p ps=0u
M1003 a_575_305# a_2463_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1004 Q_N a_575_305# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.2449e+12p ps=1.863e+07u
M1005 VPWR DE a_161_394# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 a_27_90# a_575_305# a_533_113# VNB nlowvt w=420000u l=150000u
+  ad=3.276e+11p pd=3.24e+06u as=1.008e+11p ps=1.32e+06u
M1007 a_2650_508# a_1549_74# a_2463_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=3.115e+11p ps=2.71e+06u
M1008 a_1071_462# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1009 a_1934_508# a_1351_74# a_1747_118# VPB pshort w=420000u l=180000u
+  ad=1.05e+11p pd=1.34e+06u as=1.344e+11p ps=1.48e+06u
M1010 a_1747_118# a_1549_74# a_697_113# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=4.823e+11p ps=5.11e+06u
M1011 a_1549_74# a_1351_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_119_464# D a_27_90# VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=3.52e+11p ps=3.66e+06u
M1013 VPWR a_1972_92# a_1934_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q_N a_575_305# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 VPWR a_2463_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1016 a_1351_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1017 a_533_113# a_161_394# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_697_113# SCE a_1075_125# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 VGND DE a_161_394# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1020 VPWR a_575_305# a_2650_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_157_90# D a_27_90# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1022 VGND DE a_157_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1351_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1024 a_2391_74# a_1972_92# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1025 a_2463_74# a_1549_74# a_2391_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1026 a_559_464# DE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1027 VGND a_1972_92# a_1895_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1075_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_161_394# a_119_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_90# a_575_305# a_559_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_575_305# a_2463_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1032 a_697_113# a_667_87# a_1071_462# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_697_113# a_667_87# a_27_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2463_74# a_1351_74# a_2348_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.95e+11p ps=3.59e+06u
M1035 a_1972_92# a_1747_118# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1036 a_2565_74# a_1351_74# a_2463_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1037 VGND a_575_305# a_2565_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR SCE a_667_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.208e+11p ps=1.97e+06u
M1039 a_697_113# SCE a_27_90# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1972_92# a_1747_118# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.92e+11p pd=1.88e+06u as=0p ps=0u
M1041 VGND a_2463_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1042 VGND SCE a_667_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1043 a_2348_392# a_1972_92# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1377_368# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=3.44925e+12p ps=2.926e+07u
M1001 a_141_74# D a_32_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.835e+11p ps=3.03e+06u
M1002 VPWR a_575_87# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1003 VPWR a_183_290# a_135_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1004 a_1586_74# a_1377_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.61097e+12p ps=2.285e+07u
M1005 a_32_74# a_575_87# a_527_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VPWR a_575_87# a_2675_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_2417_74# a_2013_71# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1008 a_1586_74# a_1377_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1009 a_691_113# a_661_87# a_32_74# VNB nlowvt w=420000u l=150000u
+  ad=3.885e+11p pd=4.37e+06u as=0p ps=0u
M1010 a_2489_74# a_1586_74# a_2417_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1011 a_2591_74# a_1377_368# a_2489_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 a_575_87# a_2489_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 VPWR DE a_183_290# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1014 VPWR SCE a_661_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1015 a_1784_97# a_1586_74# a_691_113# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.76e+11p ps=5.08e+06u
M1016 VPWR a_2013_71# a_1947_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1017 a_1091_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_2013_71# a_1784_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1019 a_1947_508# a_1377_368# a_1784_97# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND DE a_183_290# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1021 a_527_113# a_183_290# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_575_87# a_2591_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_575_87# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1024 a_32_74# a_575_87# a_581_462# VPB pshort w=640000u l=180000u
+  ad=3.52e+11p pd=3.66e+06u as=1.344e+11p ps=1.7e+06u
M1025 VGND a_2013_71# a_1920_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.953e+11p ps=1.77e+06u
M1026 Q a_2489_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1027 a_135_464# D a_32_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_691_113# SCE a_32_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1377_368# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1030 a_2675_508# a_1586_74# a_2489_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.115e+11p ps=2.71e+06u
M1031 a_1091_453# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1032 a_2013_71# a_1784_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1033 a_691_113# SCE a_1091_125# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2489_74# a_1377_368# a_2377_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.75e+11p ps=3.55e+06u
M1035 a_1784_97# a_1377_368# a_691_113# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1036 Q a_2489_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1037 VGND SCE a_661_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1038 a_1920_97# a_1586_74# a_1784_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_2489_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_691_113# a_661_87# a_1091_453# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_575_87# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND DE a_141_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_2377_392# a_2013_71# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_575_87# a_2489_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1045 a_581_462# DE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Q_N a_575_87# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_2489_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 VPWR a_2385_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=2.51215e+12p pd=2.218e+07u as=2.912e+11p ps=2.76e+06u
M1001 a_557_463# DE VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1002 VGND DE a_143_74# VNB nlowvt w=420000u l=150000u
+  ad=1.9208e+12p pd=1.749e+07u as=1.008e+11p ps=1.32e+06u
M1003 VGND a_2385_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 a_1492_74# a_1295_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 a_1056_455# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1006 a_1295_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1007 VGND DE a_159_404# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1008 a_505_111# a_159_404# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 a_1910_71# a_1688_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.184e+11p pd=2.2e+06u as=0p ps=0u
M1010 a_143_74# D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.982e+11p ps=3.1e+06u
M1011 a_1295_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 a_2385_74# a_1295_74# a_2277_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=7.55e+11p ps=3.51e+06u
M1013 a_547_301# a_2385_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1014 VPWR SCE a_639_85# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1015 a_27_74# a_547_301# a_557_463# VPB pshort w=640000u l=180000u
+  ad=3.456e+11p pd=3.64e+06u as=0p ps=0u
M1016 a_2313_74# a_1910_71# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1017 a_1492_74# a_1295_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1018 a_2385_74# a_1492_74# a_2313_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1019 a_669_111# SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=4.441e+11p pd=4.97e+06u as=0p ps=0u
M1020 a_669_111# a_639_85# a_1056_455# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR DE a_159_404# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1022 a_669_111# a_639_85# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=3.843e+11p pd=4.35e+06u as=0p ps=0u
M1023 a_1688_97# a_1295_74# a_669_111# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1024 a_117_464# D a_27_74# VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1025 a_2571_508# a_1492_74# a_2385_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1026 a_1688_97# a_1492_74# a_669_111# VPB pshort w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1027 a_1893_508# a_1295_74# a_1688_97# VPB pshort w=420000u l=180000u
+  ad=1.05e+11p pd=1.34e+06u as=0p ps=0u
M1028 a_669_111# SCE a_1026_125# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1029 VGND a_1910_71# a_1824_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.806e+11p ps=1.7e+06u
M1030 VPWR a_1910_71# a_1893_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1026_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1824_97# a_1492_74# a_1688_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1910_71# a_1688_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1034 a_547_301# a_2385_74# VPWR VPB pshort w=640000u l=180000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1035 a_2487_74# a_1295_74# a_2385_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1036 VGND a_547_301# a_2487_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_547_301# a_2571_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_159_404# a_117_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_27_74# a_547_301# a_505_111# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND SCE a_639_85# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1041 a_2277_392# a_1910_71# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_2660_508# a_1538_74# a_2474_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.962e+11p ps=2.72e+06u
M1001 a_2474_74# a_1538_74# a_2402_74# VNB nlowvt w=640000u l=150000u
+  ad=1.915e+11p pd=1.93e+06u as=1.344e+11p ps=1.7e+06u
M1002 a_693_113# a_663_87# a_1082_455# VPB pshort w=640000u l=180000u
+  ad=4.728e+11p pd=5.07e+06u as=1.536e+11p ps=1.76e+06u
M1003 a_1068_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.2744e+12p ps=1.998e+07u
M1004 a_1340_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VPWR DE a_180_290# VPB pshort w=640000u l=180000u
+  ad=2.92365e+12p pd=2.518e+07u as=1.792e+11p ps=1.84e+06u
M1006 VPWR SCE a_663_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1007 a_1736_97# a_1538_74# a_693_113# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1008 a_693_113# SCE a_1068_125# VNB nlowvt w=420000u l=150000u
+  ad=3.885e+11p pd=4.37e+06u as=0p ps=0u
M1009 a_548_87# a_2474_74# VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1010 Q a_2474_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1011 a_1939_508# a_1340_74# a_1736_97# VPB pshort w=420000u l=180000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1012 a_138_74# D a_40_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.982e+11p ps=3.1e+06u
M1013 a_1538_74# a_1340_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1014 a_1979_71# a_1736_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1015 VPWR a_548_87# a_2660_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_40_464# a_548_87# a_578_463# VPB pshort w=640000u l=180000u
+  ad=3.52e+11p pd=3.66e+06u as=1.344e+11p ps=1.7e+06u
M1017 Q a_2474_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1018 a_132_464# D a_40_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_693_113# SCE a_40_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1736_97# a_1340_74# a_693_113# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1021 VGND DE a_180_290# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1022 a_2360_392# a_1979_71# VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.8e+11p pd=3.56e+06u as=0p ps=0u
M1023 a_500_113# a_180_290# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1024 VPWR a_1979_71# a_1939_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_2474_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1082_455# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1872_97# a_1538_74# a_1736_97# VNB nlowvt w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=0p ps=0u
M1028 a_1979_71# a_1736_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1029 VGND a_1979_71# a_1872_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_578_463# DE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2569_74# a_1340_74# a_2474_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1032 VGND a_548_87# a_2569_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_548_87# a_2474_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1034 a_1340_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1035 a_1538_74# a_1340_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1036 a_40_464# a_548_87# a_500_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_693_113# a_663_87# a_40_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_180_290# a_132_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND DE a_138_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND SCE a_663_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1041 VGND a_2474_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_2474_74# a_1340_74# a_2360_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_2402_74# a_1979_71# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_2589_508# a_1510_74# a_2403_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.836e+11p ps=2.66e+06u
M1001 a_575_463# DE VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=3.10925e+12p ps=2.772e+07u
M1002 a_135_74# D a_37_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.373e+11p ps=2.81e+06u
M1003 a_661_113# SCE a_1044_125# VNB nlowvt w=420000u l=150000u
+  ad=5.502e+11p pd=5.14e+06u as=8.82e+10p ps=1.26e+06u
M1004 a_129_464# D a_37_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=3.52e+11p ps=3.66e+06u
M1005 a_1074_455# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1006 VGND DE a_177_290# VNB nlowvt w=420000u l=150000u
+  ad=2.3264e+12p pd=2.159e+07u as=1.197e+11p ps=1.41e+06u
M1007 a_1044_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_545_87# a_2589_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_177_290# a_129_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1313_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1011 a_1510_74# a_1313_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 Q a_2403_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1013 a_2498_74# a_1313_74# a_2403_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.915e+11p ps=1.93e+06u
M1014 VGND a_545_87# a_2498_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1510_74# a_1313_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1016 a_545_87# a_2403_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1017 Q a_2403_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=4.11e+06u as=0p ps=0u
M1018 a_37_464# a_545_87# a_497_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 a_661_113# a_631_87# a_37_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1313_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1021 a_1943_53# a_1756_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.184e+11p pd=2.2e+06u as=0p ps=0u
M1022 a_2403_74# a_1510_74# a_2331_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1023 a_37_464# a_545_87# a_575_463# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR SCE a_631_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1025 VGND a_1943_53# a_1858_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.785e+11p ps=1.69e+06u
M1026 VGND DE a_135_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_661_113# SCE a_37_464# VPB pshort w=640000u l=180000u
+  ad=4.452e+11p pd=4.97e+06u as=0p ps=0u
M1028 a_661_113# a_631_87# a_1074_455# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR DE a_177_290# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1030 a_545_87# a_2403_74# VPWR VPB pshort w=640000u l=180000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1031 a_1858_79# a_1510_74# a_1756_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.6695e+11p ps=1.74e+06u
M1032 VPWR a_2403_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1756_97# a_1510_74# a_661_113# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1034 a_497_113# a_177_290# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_2403_74# a_1313_74# a_2295_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.8e+11p ps=3.56e+06u
M1036 VPWR a_1943_53# a_1902_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1037 VGND a_2403_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1756_97# a_1313_74# a_661_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Q a_2403_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_2403_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Q a_2403_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1902_508# a_1313_74# a_1756_97# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND SCE a_631_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1044 a_2295_392# a_1943_53# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR a_2403_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1943_53# a_1756_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1047 a_2331_74# a_1943_53# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__tap_1 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__tap_2 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__tapmet1_2 VGND VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__tapvgnd_1 VGND VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__tapvgnd2_1 VGND VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__tapvpwrvgnd_1 VGND VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor2_1 A B VGND VNB VPB VPWR Y
M1000 VGND A a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=5.4e+11p pd=4.52e+06u as=4.107e+11p ps=4.07e+06u
M1001 VPWR B a_141_385# VPB pshort w=840000u l=180000u
+  ad=1.13705e+12p pd=8.5e+06u as=2.268e+11p ps=2.22e+06u
M1002 a_141_385# B a_112_119# VNB nlowvt w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=1.344e+11p ps=1.7e+06u
M1003 a_379_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1004 Y a_141_385# a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=2.294e+11p pd=2.1e+06u as=0p ps=0u
M1005 Y B a_379_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1006 a_112_119# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_141_385# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_293_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_141_385# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor2_2 A B VGND VNB VPB VPWR Y
M1000 Y B a_641_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=8.894e+11p ps=6.2e+06u
M1001 a_340_107# B VGND VNB nlowvt w=740000u l=150000u
+  ad=8.30525e+11p pd=8.22e+06u as=1.024e+12p ps=7.92e+06u
M1002 VPWR A a_641_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.16185e+12p pd=1.301e+07u as=0p ps=0u
M1003 a_641_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_136_368# a_340_107# VNB nlowvt w=740000u l=150000u
+  ad=4.008e+11p pd=2.67e+06u as=0p ps=0u
M1005 VGND B a_340_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_340_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_340_107# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_641_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_136_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_136_368# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_136_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1012 VPWR B a_136_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_136_368# B a_151_74# VNB nlowvt w=740000u l=150000u
+  ad=2.06875e+11p pd=2.05e+06u as=1.776e+11p ps=1.96e+06u
M1014 a_151_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_340_107# a_136_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor2_4 A B VGND VNB VPB VPWR Y
M1000 a_950_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.5344e+12p pd=1.394e+07u as=2.62112e+12p ps=1.87e+07u
M1001 VGND B a_511_74# VNB nlowvt w=740000u l=150000u
+  ad=1.7674e+12p pd=1.293e+07u as=1.6317e+12p ps=1.477e+07u
M1002 a_511_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B a_950_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.072e+11p pd=8.34e+06u as=0p ps=0u
M1004 a_950_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_950_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_950_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_950_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B a_950_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_511_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_511_74# a_119_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1011 a_950_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_119_368# A VPWR VPB pshort w=840000u l=180000u
+  ad=4.536e+11p pd=4.44e+06u as=0p ps=0u
M1013 VPWR A a_119_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_511_74# a_119_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_511_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_511_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_119_368# a_511_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_119_368# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# A VGND VNB nlowvt w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=0p ps=0u
M1020 VPWR B a_119_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A a_511_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_74# B a_119_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1023 a_511_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_511_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y a_119_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_119_368# B a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_119_368# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_119_368# a_511_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor3_1 A B C VGND VNB VPB VPWR X
M1000 a_81_268# C a_363_394# VPB pshort w=840000u l=180000u
+  ad=3.9275e+11p pd=2.79e+06u as=5.184e+11p ps=4.63e+06u
M1001 a_786_100# B VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.0267e+12p ps=7.95e+06u
M1002 a_786_100# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.212e+12p ps=9e+06u
M1003 VGND a_81_268# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 a_1116_383# B a_371_74# VNB nlowvt w=640000u l=150000u
+  ad=4.096e+11p pd=3.95e+06u as=4.48e+11p ps=3.96e+06u
M1005 a_1116_383# a_897_54# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_363_394# a_232_162# a_81_268# VNB nlowvt w=640000u l=150000u
+  ad=4.271e+11p pd=3.96e+06u as=2.24e+11p ps=1.98e+06u
M1007 a_371_74# a_786_100# a_897_54# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.95425e+11p ps=4.74e+06u
M1008 a_81_268# C a_371_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_363_394# a_786_100# a_897_54# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=6.9725e+11p ps=5.56e+06u
M1010 a_1116_383# B a_363_394# VPB pshort w=640000u l=180000u
+  ad=4.578e+11p pd=4.39e+06u as=0p ps=0u
M1011 a_1116_383# a_897_54# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_371_74# a_786_100# a_1116_383# VPB pshort w=640000u l=180000u
+  ad=5.792e+11p pd=4.82e+06u as=0p ps=0u
M1013 a_232_162# C VGND VNB nlowvt w=420000u l=150000u
+  ad=1.575e+11p pd=1.59e+06u as=0p ps=0u
M1014 a_897_54# B a_363_394# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_897_54# B a_371_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_81_268# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1017 VGND A a_897_54# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_232_162# C VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1019 a_371_74# a_232_162# a_81_268# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_897_54# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_363_394# a_786_100# a_1116_383# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor3_2 A B C VGND VNB VPB VPWR X
M1000 a_335_373# B a_83_247# VPB pshort w=840000u l=180000u
+  ad=5.572e+11p pd=4.77e+06u as=7.096e+11p ps=5.58e+06u
M1001 a_83_247# a_397_21# a_329_81# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=5.174e+11p ps=4.63e+06u
M1002 a_83_247# a_397_21# a_335_373# VNB nlowvt w=640000u l=150000u
+  ad=5.925e+11p pd=4.86e+06u as=4.512e+11p ps=3.97e+06u
M1003 a_335_373# B a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.886e+11p ps=3.85e+06u
M1004 a_27_373# a_397_21# a_329_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.22e+11p ps=4.25e+06u
M1005 a_1057_74# a_1027_48# a_335_373# VPB pshort w=840000u l=180000u
+  ad=4.0245e+11p pd=2.81e+06u as=0p ps=0u
M1006 X a_1057_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.5438e+12p ps=1.187e+07u
M1007 a_329_81# C a_1057_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_1057_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_1057_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.54235e+12p ps=1.041e+07u
M1010 a_83_247# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_373# a_397_21# a_335_373# VPB pshort w=640000u l=180000u
+  ad=4.656e+11p pd=4.42e+06u as=0p ps=0u
M1012 VGND a_83_247# a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C a_1027_48# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1014 a_329_81# B a_27_373# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_83_247# a_27_373# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_397_21# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 VGND a_1057_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_329_81# B a_83_247# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_335_373# C a_1057_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1020 VPWR C a_1027_48# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1021 VPWR B a_397_21# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1022 a_83_247# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1057_74# a_1027_48# a_329_81# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor3_4 A B C VGND VNB VPB VPWR X
M1000 a_75_227# a_386_23# a_321_77# VPB pshort w=840000u l=180000u
+  ad=7.2195e+11p pd=5.6e+06u as=4.964e+11p ps=4.58e+06u
M1001 X a_1057_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=2.35215e+12p ps=1.359e+07u
M1002 X a_1057_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=2.2864e+12p ps=1.53e+07u
M1003 a_75_227# A VGND VNB nlowvt w=640000u l=150000u
+  ad=5.611e+11p pd=4.74e+06u as=0p ps=0u
M1004 X a_1057_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_327_373# B a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=3.84e+11p pd=3.76e+06u as=4.635e+11p ps=4.06e+06u
M1006 a_27_373# a_386_23# a_321_77# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.739e+11p ps=3.78e+06u
M1007 VPWR B a_386_23# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 VPWR a_1057_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_75_227# a_386_23# a_327_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_327_373# C a_1057_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.592e+11p ps=2.09e+06u
M1011 VGND a_1057_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C a_1024_300# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1013 VGND a_1057_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_373# a_386_23# a_327_373# VPB pshort w=640000u l=180000u
+  ad=4.528e+11p pd=4.38e+06u as=6.18e+11p ps=4.96e+06u
M1015 a_321_77# B a_27_373# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_75_227# a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND C a_1024_300# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 a_75_227# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_321_77# C a_1057_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.305e+11p ps=2.98e+06u
M1020 VPWR a_75_227# a_27_373# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1057_74# a_1024_300# a_327_373# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B a_386_23# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 X a_1057_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_321_77# B a_75_227# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_327_373# B a_75_227# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1057_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1057_74# a_1024_300# a_321_77# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor2_1 A B VGND VNB VPB VPWR X
M1000 a_161_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=7.168e+11p ps=5.58e+06u
M1001 a_194_125# B a_161_392# VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1002 VGND B a_194_125# VNB nlowvt w=550000u l=150000u
+  ad=8.846e+11p pd=6.8e+06u as=3.5475e+11p ps=2.39e+06u
M1003 VPWR A a_355_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=7.168e+11p ps=5.76e+06u
M1004 a_455_87# A VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1005 X B a_455_87# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1006 a_355_368# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_194_125# a_355_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.696e+11p pd=2.9e+06u as=0p ps=0u
M1008 a_194_125# A VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_194_125# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor2_2 A B VGND VNB VPB VPWR X
M1000 a_313_368# a_183_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.2432e+12p pd=1.118e+07u as=3.024e+11p ps=2.78e+06u
M1001 a_119_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=9.968e+11p ps=8.32e+06u
M1002 VPWR B a_313_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_313_368# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B a_183_74# VNB nlowvt w=640000u l=150000u
+  ad=1.4793e+12p pd=8.78e+06u as=1.792e+11p ps=1.84e+06u
M1005 a_183_74# B a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1006 X B a_399_74# VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=5.66e+11p ps=4.61e+06u
M1007 a_399_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_183_74# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_399_74# B X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_399_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_183_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_313_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_313_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_183_74# a_313_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor2_4 A B VGND VNB VPB VPWR X
M1000 VPWR B a_514_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.95185e+12p pd=1.524e+07u as=2.1112e+12p ps=1.945e+07u
M1001 a_160_98# A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.958e+11p pd=4.3e+06u as=2.40945e+12p ps=1.687e+07u
M1002 a_514_368# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_514_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_36_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.1e+11p pd=7.62e+06u as=0p ps=0u
M1005 VPWR B a_514_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_514_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_160_98# B a_36_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1008 a_514_368# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_36_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X B a_877_74# VNB nlowvt w=740000u l=150000u
+  ad=8.325e+11p pd=6.69e+06u as=1.0952e+12p ps=1.036e+07u
M1011 a_36_392# B a_160_98# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_877_74# B X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_160_98# a_514_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1014 VGND a_160_98# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_877_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_877_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_514_368# a_160_98# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_160_98# a_514_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_514_368# a_160_98# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_877_74# B X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A a_514_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A a_160_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_160_98# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X B a_877_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_877_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_514_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A a_877_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND B a_160_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_160_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor3_1 A B C VGND VNB VPB VPWR X
M1000 a_84_108# A VGND VNB nlowvt w=640000u l=150000u
+  ad=6.252e+11p pd=4.99e+06u as=1.3258e+12p ps=8.35e+06u
M1001 a_1218_396# a_1157_298# a_416_86# VPB pshort w=840000u l=180000u
+  ad=4.83e+11p pd=2.83e+06u as=5.8575e+11p ps=4.8e+06u
M1002 a_84_108# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.354e+11p pd=5.57e+06u as=1.2444e+12p ps=9e+06u
M1003 a_387_392# C a_1218_396# VPB pshort w=840000u l=180000u
+  ad=5.436e+11p pd=4.69e+06u as=0p ps=0u
M1004 X a_1218_396# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 VPWR a_84_108# a_27_134# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.656e+11p ps=4.42e+06u
M1006 a_27_134# a_452_288# a_416_86# VNB nlowvt w=420000u l=150000u
+  ad=4.987e+11p pd=4.17e+06u as=4.475e+11p ps=4.01e+06u
M1007 a_416_86# C a_1218_396# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.392e+11p ps=2.34e+06u
M1008 a_27_134# a_452_288# a_387_392# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_416_86# B a_27_134# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_84_108# a_452_288# a_416_86# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_452_288# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.035e+11p ps=2.03e+06u
M1012 a_387_392# B a_84_108# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR C a_1157_298# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.432e+11p ps=2.04e+06u
M1014 a_387_392# B a_27_134# VNB nlowvt w=640000u l=150000u
+  ad=5.1415e+11p pd=4.38e+06u as=0p ps=0u
M1015 a_416_86# B a_84_108# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1218_396# a_1157_298# a_387_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND C a_1157_298# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 X a_1218_396# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 VGND a_84_108# a_27_134# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_84_108# a_452_288# a_387_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR B a_452_288# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor3_2 A B C VGND VNB VPB VPWR X
M1000 a_83_289# A VGND VNB nlowvt w=640000u l=150000u
+  ad=6.24525e+11p pd=4.72e+06u as=1.66725e+12p ps=1.089e+07u
M1001 a_27_134# a_440_315# a_375_419# VPB pshort w=640000u l=180000u
+  ad=4.528e+11p pd=4.38e+06u as=4.932e+11p ps=4.57e+06u
M1002 VGND a_1198_424# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1003 a_416_113# B a_27_134# VPB pshort w=640000u l=180000u
+  ad=5.184e+11p pd=4.63e+06u as=0p ps=0u
M1004 X a_1198_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.807e+12p ps=1.21e+07u
M1005 a_1198_424# a_1162_379# a_375_419# VNB nlowvt w=640000u l=150000u
+  ad=3.3955e+11p pd=2.48e+06u as=4.75e+11p ps=4.11e+06u
M1006 VPWR a_83_289# a_27_134# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_1198_424# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_83_289# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.848e+11p pd=5.68e+06u as=0p ps=0u
M1009 a_416_113# C a_1198_424# VNB nlowvt w=640000u l=150000u
+  ad=4.219e+11p pd=3.93e+06u as=0p ps=0u
M1010 a_27_134# a_440_315# a_416_113# VNB nlowvt w=420000u l=150000u
+  ad=4.987e+11p pd=4.17e+06u as=0p ps=0u
M1011 VGND B a_440_315# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.035e+11p ps=2.03e+06u
M1012 a_375_419# C a_1198_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.872e+11p ps=2.84e+06u
M1013 a_83_289# a_440_315# a_416_113# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_1198_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1198_424# a_1162_379# a_416_113# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR C a_1162_379# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.304e+11p ps=2e+06u
M1017 a_375_419# B a_27_134# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_83_289# a_27_134# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C a_1162_379# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1020 a_416_113# B a_83_289# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_83_289# a_440_315# a_375_419# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR B a_440_315# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1023 a_375_419# B a_83_289# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor3_4 A B C VGND VNB VPB VPWR X
M1000 VPWR C a_1155_284# VPB pshort w=640000u l=180000u
+  ad=2.1152e+12p pd=1.487e+07u as=1.792e+11p ps=1.84e+06u
M1001 VGND C a_1155_284# VNB nlowvt w=420000u l=150000u
+  ad=1.6131e+12p pd=1.223e+07u as=2.121e+11p ps=1.85e+06u
M1002 VPWR a_74_294# a_27_118# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6055e+11p ps=4.93e+06u
M1003 a_1221_388# a_1155_284# a_416_118# VPB pshort w=840000u l=180000u
+  ad=4.2e+11p pd=2.68e+06u as=6.5265e+11p ps=4.95e+06u
M1004 VGND a_1221_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1005 VGND a_74_294# a_27_118# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.264e+11p ps=4.03e+06u
M1006 a_326_392# B a_27_118# VNB nlowvt w=640000u l=150000u
+  ad=4.6775e+11p pd=4.06e+06u as=0p ps=0u
M1007 a_326_392# C a_1221_388# VPB pshort w=840000u l=180000u
+  ad=5.184e+11p pd=4.63e+06u as=0p ps=0u
M1008 a_1221_388# a_1155_284# a_326_392# VNB nlowvt w=640000u l=150000u
+  ad=3.392e+11p pd=2.34e+06u as=0p ps=0u
M1009 a_326_392# B a_74_294# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=8.764e+11p ps=5.66e+06u
M1010 X a_1221_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_1221_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_1221_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1013 a_416_118# B a_74_294# VNB nlowvt w=640000u l=150000u
+  ad=3.899e+11p pd=3.83e+06u as=7.264e+11p ps=4.83e+06u
M1014 a_74_294# a_397_320# a_416_118# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B a_397_320# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1016 a_416_118# C a_1221_388# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_1221_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_118# a_397_320# a_416_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_118# a_397_320# a_326_392# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1221_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_416_118# B a_27_118# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1221_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_74_294# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B a_397_320# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1025 a_74_294# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1221_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_74_294# a_397_320# a_326_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0




******* EOF

