magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 920 561
rect 139 442 216 527
rect 17 199 115 340
rect 422 442 499 527
rect 705 442 782 527
rect 816 299 903 493
rect 831 165 903 299
rect 139 17 216 97
rect 422 17 499 97
rect 705 17 782 97
rect 816 51 903 165
rect 0 -17 920 17
<< obsli1 >>
rect 17 408 105 493
rect 17 374 216 408
rect 149 265 216 374
rect 250 335 304 493
rect 338 408 388 493
rect 338 369 499 408
rect 250 299 395 335
rect 149 199 231 265
rect 265 199 395 299
rect 429 265 499 369
rect 533 335 583 493
rect 617 408 671 493
rect 617 369 782 408
rect 533 299 678 335
rect 429 199 514 265
rect 548 199 678 299
rect 712 265 782 369
rect 712 199 797 265
rect 149 165 216 199
rect 265 165 304 199
rect 429 165 499 199
rect 548 165 583 199
rect 712 165 782 199
rect 17 131 216 165
rect 17 51 105 131
rect 250 51 304 165
rect 338 131 499 165
rect 338 51 388 131
rect 533 51 583 165
rect 617 131 782 165
rect 617 51 671 131
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 17 199 115 340 6 A
port 1 nsew signal input
rlabel locali s 831 165 903 299 6 X
port 2 nsew signal output
rlabel locali s 816 299 903 493 6 X
port 2 nsew signal output
rlabel locali s 816 51 903 165 6 X
port 2 nsew signal output
rlabel locali s 705 17 782 97 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 422 17 499 97 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 139 17 216 97 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 920 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 705 442 782 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 422 442 499 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 139 442 216 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 920 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 920 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2846780
string GDS_START 2839256
<< end >>
