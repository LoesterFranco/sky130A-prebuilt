magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 25 236 75 596
rect 109 270 175 356
rect 217 270 359 356
rect 393 270 459 356
rect 501 270 567 356
rect 601 236 743 310
rect 25 202 515 236
rect 25 70 218 202
rect 432 70 515 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 115 581 411 615
rect 115 390 181 581
rect 255 424 309 547
rect 345 458 411 581
rect 451 424 501 596
rect 535 458 605 649
rect 639 424 705 596
rect 255 390 705 424
rect 639 364 705 390
rect 252 17 326 165
rect 634 17 700 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 501 270 567 356 6 A1
port 1 nsew signal input
rlabel locali s 601 236 743 310 6 A2
port 2 nsew signal input
rlabel locali s 393 270 459 356 6 B1
port 3 nsew signal input
rlabel locali s 217 270 359 356 6 B2
port 4 nsew signal input
rlabel locali s 109 270 175 356 6 C1
port 5 nsew signal input
rlabel locali s 432 70 515 202 6 Y
port 6 nsew signal output
rlabel locali s 25 236 75 596 6 Y
port 6 nsew signal output
rlabel locali s 25 202 515 236 6 Y
port 6 nsew signal output
rlabel locali s 25 70 218 202 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3535912
string GDS_START 3528054
<< end >>
