magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 51 367 102 527
rect 136 333 202 493
rect 236 367 270 527
rect 304 333 370 493
rect 404 367 438 527
rect 472 333 538 493
rect 572 367 606 527
rect 640 333 706 493
rect 740 367 800 527
rect 17 299 811 333
rect 17 181 86 299
rect 136 215 707 265
rect 747 181 811 299
rect 17 143 811 181
rect 51 17 102 109
rect 136 51 202 143
rect 236 17 270 109
rect 304 51 370 143
rect 404 17 438 109
rect 472 51 538 143
rect 572 17 606 109
rect 640 51 706 143
rect 740 17 801 109
rect 0 -17 828 17
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 136 215 707 265 6 A
port 1 nsew signal input
rlabel locali s 747 181 811 299 6 Y
port 2 nsew signal output
rlabel locali s 640 333 706 493 6 Y
port 2 nsew signal output
rlabel locali s 640 51 706 143 6 Y
port 2 nsew signal output
rlabel locali s 472 333 538 493 6 Y
port 2 nsew signal output
rlabel locali s 472 51 538 143 6 Y
port 2 nsew signal output
rlabel locali s 304 333 370 493 6 Y
port 2 nsew signal output
rlabel locali s 304 51 370 143 6 Y
port 2 nsew signal output
rlabel locali s 136 333 202 493 6 Y
port 2 nsew signal output
rlabel locali s 136 51 202 143 6 Y
port 2 nsew signal output
rlabel locali s 17 299 811 333 6 Y
port 2 nsew signal output
rlabel locali s 17 181 86 299 6 Y
port 2 nsew signal output
rlabel locali s 17 143 811 181 6 Y
port 2 nsew signal output
rlabel locali s 740 17 801 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 572 17 606 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 404 17 438 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 236 17 270 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 51 17 102 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 740 367 800 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 572 367 606 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 404 367 438 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 236 367 270 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 51 367 102 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2224192
string GDS_START 2216692
<< end >>
