magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1288 561
rect 35 289 69 527
rect 307 357 341 527
rect 475 357 509 527
rect 543 323 609 493
rect 643 367 677 527
rect 711 323 777 493
rect 811 367 845 527
rect 879 323 945 493
rect 979 367 1013 527
rect 1047 323 1113 493
rect 1147 367 1181 527
rect 543 289 1271 323
rect 17 215 101 255
rect 1194 181 1271 289
rect 35 17 69 181
rect 543 147 1271 181
rect 307 17 341 113
rect 475 17 509 113
rect 543 52 609 147
rect 643 17 677 113
rect 711 52 777 147
rect 811 17 845 113
rect 879 52 945 147
rect 979 17 1013 113
rect 1047 52 1113 147
rect 1147 17 1181 113
rect 0 -17 1288 17
<< obsli1 >>
rect 103 309 169 493
rect 135 255 169 309
rect 207 323 273 493
rect 375 323 441 493
rect 207 289 509 323
rect 475 255 509 289
rect 135 215 441 255
rect 475 215 1152 255
rect 135 181 169 215
rect 475 181 509 215
rect 103 52 169 181
rect 207 147 509 181
rect 207 52 273 147
rect 375 52 441 147
<< metal1 >>
rect 0 496 1288 592
rect 0 -48 1288 48
<< labels >>
rlabel locali s 17 215 101 255 6 A
port 1 nsew signal input
rlabel locali s 1194 181 1271 289 6 Y
port 2 nsew signal output
rlabel locali s 1047 323 1113 493 6 Y
port 2 nsew signal output
rlabel locali s 1047 52 1113 147 6 Y
port 2 nsew signal output
rlabel locali s 879 323 945 493 6 Y
port 2 nsew signal output
rlabel locali s 879 52 945 147 6 Y
port 2 nsew signal output
rlabel locali s 711 323 777 493 6 Y
port 2 nsew signal output
rlabel locali s 711 52 777 147 6 Y
port 2 nsew signal output
rlabel locali s 543 323 609 493 6 Y
port 2 nsew signal output
rlabel locali s 543 289 1271 323 6 Y
port 2 nsew signal output
rlabel locali s 543 147 1271 181 6 Y
port 2 nsew signal output
rlabel locali s 543 52 609 147 6 Y
port 2 nsew signal output
rlabel locali s 1147 17 1181 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 979 17 1013 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 811 17 845 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 643 17 677 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 475 17 509 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 307 17 341 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 35 17 69 181 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1288 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1147 367 1181 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 979 367 1013 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 811 367 845 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 643 367 677 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 475 357 509 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 307 357 341 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 35 289 69 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 1288 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3113144
string GDS_START 3102992
<< end >>
