magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 2630 704
rect 193 322 1347 332
rect 1139 305 1347 322
<< pwell >>
rect 0 0 2592 49
<< scpmos >>
rect 86 508 116 592
rect 288 358 318 582
rect 378 358 408 582
rect 586 463 616 547
rect 676 463 706 547
rect 760 463 790 547
rect 945 463 975 547
rect 1048 463 1078 547
rect 1228 341 1258 541
rect 1329 392 1359 592
rect 1491 508 1521 592
rect 1575 508 1605 592
rect 1665 508 1695 592
rect 1882 368 1912 452
rect 1989 368 2019 592
rect 2079 368 2109 592
rect 2280 368 2310 568
rect 2386 368 2416 592
rect 2476 368 2506 592
<< nmoslvt >>
rect 84 74 114 158
rect 282 74 312 222
rect 368 74 398 222
rect 565 97 595 181
rect 701 97 731 181
rect 773 97 803 181
rect 971 74 1001 158
rect 1043 74 1073 158
rect 1231 74 1261 202
rect 1309 74 1339 202
rect 1423 118 1453 202
rect 1501 118 1531 202
rect 1579 118 1609 202
rect 1780 118 1810 202
rect 1994 74 2024 222
rect 2080 74 2110 222
rect 2278 74 2308 202
rect 2392 74 2422 222
rect 2478 74 2508 222
<< ndiff >>
rect 225 195 282 222
rect 225 161 237 195
rect 271 161 282 195
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 171 158
rect 114 99 125 133
rect 159 99 171 133
rect 114 74 171 99
rect 225 120 282 161
rect 225 86 237 120
rect 271 86 282 120
rect 225 74 282 86
rect 312 186 368 222
rect 312 152 323 186
rect 357 152 368 186
rect 312 118 368 152
rect 312 84 323 118
rect 357 84 368 118
rect 312 74 368 84
rect 398 210 454 222
rect 398 176 409 210
rect 443 176 454 210
rect 398 120 454 176
rect 398 86 409 120
rect 443 86 454 120
rect 508 169 565 181
rect 508 135 520 169
rect 554 135 565 169
rect 508 97 565 135
rect 595 156 701 181
rect 595 122 656 156
rect 690 122 701 156
rect 595 97 701 122
rect 731 97 773 181
rect 803 148 860 181
rect 1181 158 1231 202
rect 803 114 814 148
rect 848 114 860 148
rect 803 97 860 114
rect 914 133 971 158
rect 914 99 926 133
rect 960 99 971 133
rect 398 74 454 86
rect 914 74 971 99
rect 1001 74 1043 158
rect 1073 120 1231 158
rect 1073 86 1084 120
rect 1118 86 1182 120
rect 1216 86 1231 120
rect 1073 74 1231 86
rect 1261 74 1309 202
rect 1339 174 1423 202
rect 1339 140 1364 174
rect 1398 140 1423 174
rect 1339 118 1423 140
rect 1453 118 1501 202
rect 1531 118 1579 202
rect 1609 118 1780 202
rect 1810 177 1883 202
rect 1810 143 1837 177
rect 1871 143 1883 177
rect 1810 118 1883 143
rect 1937 152 1994 222
rect 1937 118 1949 152
rect 1983 118 1994 152
rect 1339 74 1389 118
rect 1624 84 1636 118
rect 1670 84 1719 118
rect 1753 84 1765 118
rect 1624 72 1765 84
rect 1937 74 1994 118
rect 2024 210 2080 222
rect 2024 176 2035 210
rect 2069 176 2080 210
rect 2024 120 2080 176
rect 2024 86 2035 120
rect 2069 86 2080 120
rect 2024 74 2080 86
rect 2110 210 2167 222
rect 2110 176 2121 210
rect 2155 176 2167 210
rect 2342 202 2392 222
rect 2110 120 2167 176
rect 2110 86 2121 120
rect 2155 86 2167 120
rect 2110 74 2167 86
rect 2221 190 2278 202
rect 2221 156 2233 190
rect 2267 156 2278 190
rect 2221 120 2278 156
rect 2221 86 2233 120
rect 2267 86 2278 120
rect 2221 74 2278 86
rect 2308 190 2392 202
rect 2308 156 2333 190
rect 2367 156 2392 190
rect 2308 120 2392 156
rect 2308 86 2333 120
rect 2367 86 2392 120
rect 2308 74 2392 86
rect 2422 210 2478 222
rect 2422 176 2433 210
rect 2467 176 2478 210
rect 2422 120 2478 176
rect 2422 86 2433 120
rect 2467 86 2478 120
rect 2422 74 2478 86
rect 2508 210 2565 222
rect 2508 176 2519 210
rect 2553 176 2565 210
rect 2508 120 2565 176
rect 2508 86 2519 120
rect 2553 86 2565 120
rect 2508 74 2565 86
<< pdiff >>
rect 27 567 86 592
rect 27 533 39 567
rect 73 533 86 567
rect 27 508 86 533
rect 116 568 175 592
rect 116 534 129 568
rect 163 534 175 568
rect 116 508 175 534
rect 229 404 288 582
rect 229 370 241 404
rect 275 370 288 404
rect 229 358 288 370
rect 318 563 378 582
rect 318 529 331 563
rect 365 529 378 563
rect 318 358 378 529
rect 408 550 467 582
rect 408 516 421 550
rect 455 516 467 550
rect 408 358 467 516
rect 808 581 866 593
rect 808 547 820 581
rect 854 547 866 581
rect 1144 556 1210 568
rect 1144 547 1160 556
rect 527 520 586 547
rect 527 486 539 520
rect 573 486 586 520
rect 527 463 586 486
rect 616 520 676 547
rect 616 486 629 520
rect 663 486 676 520
rect 616 463 676 486
rect 706 463 760 547
rect 790 463 945 547
rect 975 520 1048 547
rect 975 486 988 520
rect 1022 486 1048 520
rect 975 463 1048 486
rect 1078 522 1160 547
rect 1194 541 1210 556
rect 1276 541 1329 592
rect 1194 522 1228 541
rect 1078 463 1228 522
rect 1175 341 1228 463
rect 1258 392 1329 541
rect 1359 580 1491 592
rect 1359 546 1372 580
rect 1406 546 1444 580
rect 1478 546 1491 580
rect 1359 512 1491 546
rect 1359 478 1372 512
rect 1406 508 1491 512
rect 1521 508 1575 592
rect 1605 580 1665 592
rect 1605 546 1618 580
rect 1652 546 1665 580
rect 1605 508 1665 546
rect 1695 567 1753 592
rect 1695 533 1708 567
rect 1742 533 1753 567
rect 1695 508 1753 533
rect 1930 578 1989 592
rect 1930 544 1942 578
rect 1976 544 1989 578
rect 1807 508 1864 520
rect 1406 478 1418 508
rect 1359 444 1418 478
rect 1359 410 1372 444
rect 1406 410 1418 444
rect 1359 392 1418 410
rect 1258 341 1311 392
rect 1807 474 1819 508
rect 1853 474 1864 508
rect 1807 452 1864 474
rect 1930 452 1989 544
rect 1807 368 1882 452
rect 1912 368 1989 452
rect 2019 578 2079 592
rect 2019 544 2032 578
rect 2066 544 2079 578
rect 2019 496 2079 544
rect 2019 462 2032 496
rect 2066 462 2079 496
rect 2019 414 2079 462
rect 2019 380 2032 414
rect 2066 380 2079 414
rect 2019 368 2079 380
rect 2109 578 2167 592
rect 2109 544 2122 578
rect 2156 544 2167 578
rect 2328 568 2386 592
rect 2109 496 2167 544
rect 2109 462 2122 496
rect 2156 462 2167 496
rect 2109 414 2167 462
rect 2109 380 2122 414
rect 2156 380 2167 414
rect 2109 368 2167 380
rect 2221 556 2280 568
rect 2221 522 2233 556
rect 2267 522 2280 556
rect 2221 485 2280 522
rect 2221 451 2233 485
rect 2267 451 2280 485
rect 2221 414 2280 451
rect 2221 380 2233 414
rect 2267 380 2280 414
rect 2221 368 2280 380
rect 2310 556 2386 568
rect 2310 522 2339 556
rect 2373 522 2386 556
rect 2310 485 2386 522
rect 2310 451 2339 485
rect 2373 451 2386 485
rect 2310 414 2386 451
rect 2310 380 2339 414
rect 2373 380 2386 414
rect 2310 368 2386 380
rect 2416 580 2476 592
rect 2416 546 2429 580
rect 2463 546 2476 580
rect 2416 497 2476 546
rect 2416 463 2429 497
rect 2463 463 2476 497
rect 2416 414 2476 463
rect 2416 380 2429 414
rect 2463 380 2476 414
rect 2416 368 2476 380
rect 2506 580 2565 592
rect 2506 546 2519 580
rect 2553 546 2565 580
rect 2506 497 2565 546
rect 2506 463 2519 497
rect 2553 463 2565 497
rect 2506 414 2565 463
rect 2506 380 2519 414
rect 2553 380 2565 414
rect 2506 368 2565 380
<< ndiffc >>
rect 237 161 271 195
rect 39 99 73 133
rect 125 99 159 133
rect 237 86 271 120
rect 323 152 357 186
rect 323 84 357 118
rect 409 176 443 210
rect 409 86 443 120
rect 520 135 554 169
rect 656 122 690 156
rect 814 114 848 148
rect 926 99 960 133
rect 1084 86 1118 120
rect 1182 86 1216 120
rect 1364 140 1398 174
rect 1837 143 1871 177
rect 1949 118 1983 152
rect 1636 84 1670 118
rect 1719 84 1753 118
rect 2035 176 2069 210
rect 2035 86 2069 120
rect 2121 176 2155 210
rect 2121 86 2155 120
rect 2233 156 2267 190
rect 2233 86 2267 120
rect 2333 156 2367 190
rect 2333 86 2367 120
rect 2433 176 2467 210
rect 2433 86 2467 120
rect 2519 176 2553 210
rect 2519 86 2553 120
<< pdiffc >>
rect 39 533 73 567
rect 129 534 163 568
rect 241 370 275 404
rect 331 529 365 563
rect 421 516 455 550
rect 820 547 854 581
rect 539 486 573 520
rect 629 486 663 520
rect 988 486 1022 520
rect 1160 522 1194 556
rect 1372 546 1406 580
rect 1444 546 1478 580
rect 1372 478 1406 512
rect 1618 546 1652 580
rect 1708 533 1742 567
rect 1942 544 1976 578
rect 1372 410 1406 444
rect 1819 474 1853 508
rect 2032 544 2066 578
rect 2032 462 2066 496
rect 2032 380 2066 414
rect 2122 544 2156 578
rect 2122 462 2156 496
rect 2122 380 2156 414
rect 2233 522 2267 556
rect 2233 451 2267 485
rect 2233 380 2267 414
rect 2339 522 2373 556
rect 2339 451 2373 485
rect 2339 380 2373 414
rect 2429 546 2463 580
rect 2429 463 2463 497
rect 2429 380 2463 414
rect 2519 546 2553 580
rect 2519 463 2553 497
rect 2519 380 2553 414
<< poly >>
rect 86 592 116 618
rect 482 615 1362 645
rect 288 582 318 608
rect 378 582 408 608
rect 86 493 116 508
rect 83 398 119 493
rect 83 382 161 398
rect 83 348 111 382
rect 145 348 161 382
rect 83 314 161 348
rect 288 343 318 358
rect 378 343 408 358
rect 83 280 111 314
rect 145 280 161 314
rect 285 310 321 343
rect 375 326 411 343
rect 482 326 512 615
rect 586 547 616 573
rect 673 562 709 615
rect 1326 607 1362 615
rect 1329 592 1359 607
rect 1491 592 1521 618
rect 1575 592 1605 618
rect 1665 592 1695 618
rect 1989 592 2019 618
rect 2079 592 2109 618
rect 676 547 706 562
rect 760 547 790 573
rect 945 547 975 573
rect 1048 547 1078 573
rect 1228 541 1258 567
rect 586 448 616 463
rect 583 421 619 448
rect 676 437 706 463
rect 760 448 790 463
rect 945 448 975 463
rect 1048 448 1078 463
rect 757 431 793 448
rect 368 310 512 326
rect 83 246 161 280
rect 83 212 111 246
rect 145 212 161 246
rect 260 294 326 310
rect 260 260 276 294
rect 310 260 326 294
rect 260 244 326 260
rect 368 276 405 310
rect 439 276 512 310
rect 557 405 623 421
rect 557 371 573 405
rect 607 371 623 405
rect 757 415 894 431
rect 757 401 844 415
rect 557 353 623 371
rect 828 381 844 401
rect 878 381 894 415
rect 828 365 894 381
rect 942 377 978 448
rect 1045 404 1081 448
rect 1045 388 1111 404
rect 557 337 780 353
rect 557 303 573 337
rect 607 303 730 337
rect 764 303 780 337
rect 557 287 780 303
rect 368 260 512 276
rect 282 222 312 244
rect 368 222 398 260
rect 482 239 512 260
rect 83 196 161 212
rect 84 158 114 196
rect 482 209 595 239
rect 565 181 595 209
rect 701 181 731 287
rect 859 269 889 365
rect 937 361 1003 377
rect 937 327 953 361
rect 987 327 1003 361
rect 937 311 1003 327
rect 1045 354 1061 388
rect 1095 354 1111 388
rect 1045 338 1111 354
rect 1491 493 1521 508
rect 1575 493 1605 508
rect 1665 493 1695 508
rect 1488 470 1524 493
rect 1450 454 1524 470
rect 1450 420 1466 454
rect 1500 420 1524 454
rect 1450 404 1524 420
rect 1329 377 1359 392
rect 1326 362 1362 377
rect 859 253 926 269
rect 859 233 876 253
rect 773 219 876 233
rect 910 219 926 253
rect 773 203 926 219
rect 773 181 803 203
rect 971 158 1001 311
rect 1045 203 1075 338
rect 1228 326 1258 341
rect 1326 332 1453 362
rect 1572 356 1608 493
rect 1117 274 1183 290
rect 1117 240 1133 274
rect 1167 254 1183 274
rect 1225 254 1261 326
rect 1167 240 1261 254
rect 1117 224 1261 240
rect 1043 173 1075 203
rect 1231 202 1261 224
rect 1309 274 1375 290
rect 1309 240 1325 274
rect 1359 240 1375 274
rect 1309 224 1375 240
rect 1309 202 1339 224
rect 1423 202 1453 332
rect 1545 340 1611 356
rect 1545 320 1561 340
rect 1501 306 1561 320
rect 1595 306 1611 340
rect 1501 290 1611 306
rect 1662 302 1698 493
rect 1882 452 1912 478
rect 2280 568 2310 594
rect 2386 592 2416 618
rect 2476 592 2506 618
rect 1882 353 1912 368
rect 1989 353 2019 368
rect 2079 353 2109 368
rect 2280 353 2310 368
rect 2386 353 2416 368
rect 2476 353 2506 368
rect 1879 336 1915 353
rect 1780 326 1915 336
rect 1986 326 2022 353
rect 2076 326 2112 353
rect 2277 326 2313 353
rect 2383 326 2419 353
rect 2473 326 2509 353
rect 1780 320 2313 326
rect 1501 202 1531 290
rect 1662 286 1728 302
rect 1662 252 1678 286
rect 1712 252 1728 286
rect 1662 248 1728 252
rect 1579 218 1728 248
rect 1780 286 1796 320
rect 1830 286 1864 320
rect 1898 286 2313 320
rect 1780 270 2313 286
rect 2355 310 2509 326
rect 2355 276 2371 310
rect 2405 276 2509 310
rect 1579 202 1609 218
rect 1780 202 1810 270
rect 1994 222 2024 270
rect 2080 222 2110 270
rect 1043 158 1073 173
rect 84 48 114 74
rect 282 48 312 74
rect 368 48 398 74
rect 565 71 595 97
rect 701 71 731 97
rect 773 71 803 97
rect 1423 92 1453 118
rect 1501 92 1531 118
rect 1579 92 1609 118
rect 1780 92 1810 118
rect 971 48 1001 74
rect 1043 48 1073 74
rect 1231 48 1261 74
rect 1309 48 1339 74
rect 2278 202 2308 270
rect 2355 260 2509 276
rect 2392 222 2422 260
rect 2478 222 2508 260
rect 1994 48 2024 74
rect 2080 48 2110 74
rect 2278 48 2308 74
rect 2392 48 2422 74
rect 2478 48 2508 74
<< polycont >>
rect 111 348 145 382
rect 111 280 145 314
rect 111 212 145 246
rect 276 260 310 294
rect 405 276 439 310
rect 573 371 607 405
rect 844 381 878 415
rect 573 303 607 337
rect 730 303 764 337
rect 953 327 987 361
rect 1061 354 1095 388
rect 1466 420 1500 454
rect 876 219 910 253
rect 1133 240 1167 274
rect 1325 240 1359 274
rect 1561 306 1595 340
rect 1678 252 1712 286
rect 1796 286 1830 320
rect 1864 286 1898 320
rect 2371 276 2405 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 23 567 73 596
rect 23 533 39 567
rect 23 472 73 533
rect 113 568 179 649
rect 113 534 129 568
rect 163 534 179 568
rect 113 506 179 534
rect 315 563 381 649
rect 315 529 331 563
rect 365 529 381 563
rect 315 506 381 529
rect 421 581 769 615
rect 421 550 455 581
rect 421 480 455 516
rect 489 520 573 547
rect 489 486 539 520
rect 23 446 359 472
rect 489 459 573 486
rect 613 520 691 547
rect 613 486 629 520
rect 663 486 691 520
rect 613 459 691 486
rect 489 446 523 459
rect 23 438 523 446
rect 23 162 57 438
rect 325 412 523 438
rect 95 382 161 398
rect 95 348 111 382
rect 145 348 161 382
rect 95 314 161 348
rect 95 280 111 314
rect 145 280 161 314
rect 95 246 161 280
rect 95 212 111 246
rect 145 212 161 246
rect 95 196 161 212
rect 195 370 241 404
rect 275 378 291 404
rect 275 370 455 378
rect 195 344 455 370
rect 195 202 229 344
rect 389 310 455 344
rect 263 294 355 310
rect 263 260 276 294
rect 310 260 355 294
rect 389 276 405 310
rect 439 276 455 310
rect 389 260 455 276
rect 263 236 355 260
rect 409 210 443 226
rect 195 195 287 202
rect 23 133 73 162
rect 23 99 39 133
rect 23 70 73 99
rect 109 133 159 162
rect 109 99 125 133
rect 109 17 159 99
rect 195 161 237 195
rect 271 161 287 195
rect 195 120 287 161
rect 195 86 237 120
rect 271 86 287 120
rect 195 70 287 86
rect 321 186 373 202
rect 321 152 323 186
rect 357 152 373 186
rect 321 118 373 152
rect 321 84 323 118
rect 357 84 373 118
rect 321 17 373 84
rect 409 120 443 176
rect 489 185 523 412
rect 557 405 623 421
rect 557 371 573 405
rect 607 371 623 405
rect 557 337 623 371
rect 557 303 573 337
rect 607 303 623 337
rect 557 287 623 303
rect 489 169 554 185
rect 489 135 520 169
rect 489 119 554 135
rect 409 85 443 86
rect 588 85 622 287
rect 657 253 691 459
rect 725 513 769 581
rect 804 581 870 649
rect 804 547 820 581
rect 854 547 870 581
rect 904 581 1106 615
rect 904 513 938 581
rect 725 479 938 513
rect 972 520 1038 547
rect 972 486 988 520
rect 1022 486 1038 520
rect 725 337 769 479
rect 972 459 1038 486
rect 1072 472 1106 581
rect 1140 556 1214 649
rect 1140 522 1160 556
rect 1194 522 1214 556
rect 1140 506 1214 522
rect 1356 580 1494 596
rect 1356 546 1372 580
rect 1406 546 1444 580
rect 1478 546 1494 580
rect 1356 530 1494 546
rect 1618 580 1652 649
rect 1618 530 1652 546
rect 1692 567 1758 583
rect 1692 533 1708 567
rect 1742 533 1758 567
rect 1356 512 1584 530
rect 1356 478 1372 512
rect 1406 496 1584 512
rect 1692 496 1758 533
rect 1926 578 1992 649
rect 1926 544 1942 578
rect 1976 544 1992 578
rect 1926 526 1992 544
rect 2026 578 2087 594
rect 2026 544 2032 578
rect 2066 544 2087 578
rect 972 445 1006 459
rect 828 415 1006 445
rect 1072 438 1300 472
rect 828 381 844 415
rect 878 411 1006 415
rect 878 381 894 411
rect 828 371 894 381
rect 1045 388 1127 404
rect 950 361 1003 377
rect 950 337 953 361
rect 725 303 730 337
rect 764 303 769 337
rect 725 287 769 303
rect 803 327 953 337
rect 987 327 1003 361
rect 803 303 1003 327
rect 1045 354 1061 388
rect 1095 354 1127 388
rect 1045 350 1127 354
rect 1045 316 1087 350
rect 1121 316 1127 350
rect 803 253 837 303
rect 950 282 1003 303
rect 1266 290 1300 438
rect 1356 444 1406 478
rect 1356 410 1372 444
rect 1356 370 1406 410
rect 1450 454 1516 462
rect 1450 420 1466 454
rect 1500 420 1516 454
rect 1450 404 1516 420
rect 1550 424 1758 496
rect 1803 508 1869 524
rect 1803 474 1819 508
rect 1853 492 1869 508
rect 2026 496 2087 544
rect 1853 474 1982 492
rect 1803 458 1982 474
rect 1356 336 1443 370
rect 950 274 1183 282
rect 657 219 837 253
rect 871 253 916 269
rect 871 219 876 253
rect 910 219 916 253
rect 950 248 1133 274
rect 1117 240 1133 248
rect 1167 240 1183 274
rect 1117 224 1183 240
rect 1266 274 1375 290
rect 1266 240 1325 274
rect 1359 240 1375 274
rect 1266 224 1375 240
rect 657 185 706 219
rect 871 203 916 219
rect 656 156 706 185
rect 690 122 706 156
rect 656 93 706 122
rect 798 148 848 169
rect 798 114 814 148
rect 409 51 622 85
rect 798 17 848 114
rect 882 133 976 203
rect 882 99 926 133
rect 960 99 976 133
rect 882 70 976 99
rect 1068 120 1232 136
rect 1068 86 1084 120
rect 1118 86 1182 120
rect 1216 86 1232 120
rect 1068 17 1232 86
rect 1266 90 1300 224
rect 1409 190 1443 336
rect 1334 174 1443 190
rect 1334 140 1364 174
rect 1398 140 1443 174
rect 1334 124 1443 140
rect 1477 90 1511 404
rect 1550 390 1914 424
rect 1545 340 1611 356
rect 1545 306 1561 340
rect 1595 306 1611 340
rect 1545 202 1611 306
rect 1657 350 1728 356
rect 1657 316 1663 350
rect 1697 316 1728 350
rect 1657 286 1728 316
rect 1657 252 1678 286
rect 1712 252 1728 286
rect 1780 320 1914 390
rect 1780 286 1796 320
rect 1830 286 1864 320
rect 1898 286 1914 320
rect 1780 270 1914 286
rect 1657 236 1728 252
rect 1948 236 1982 458
rect 2026 462 2032 496
rect 2066 462 2087 496
rect 2026 414 2087 462
rect 2026 380 2032 414
rect 2066 380 2087 414
rect 2026 364 2087 380
rect 2121 578 2172 649
rect 2121 544 2122 578
rect 2156 544 2172 578
rect 2121 496 2172 544
rect 2121 462 2122 496
rect 2156 462 2172 496
rect 2121 414 2172 462
rect 2121 380 2122 414
rect 2156 380 2172 414
rect 2121 364 2172 380
rect 2217 556 2283 572
rect 2217 522 2233 556
rect 2267 522 2283 556
rect 2217 485 2283 522
rect 2217 451 2233 485
rect 2267 451 2283 485
rect 2217 414 2283 451
rect 2217 380 2233 414
rect 2267 380 2283 414
rect 1821 202 1982 236
rect 2035 210 2087 364
rect 2217 326 2283 380
rect 2323 556 2373 649
rect 2323 522 2339 556
rect 2323 485 2373 522
rect 2323 451 2339 485
rect 2323 414 2373 451
rect 2323 380 2339 414
rect 2323 364 2373 380
rect 2413 580 2485 596
rect 2413 546 2429 580
rect 2463 546 2485 580
rect 2413 497 2485 546
rect 2413 463 2429 497
rect 2463 463 2485 497
rect 2413 414 2485 463
rect 2413 380 2429 414
rect 2463 380 2485 414
rect 2413 364 2485 380
rect 2519 580 2569 649
rect 2553 546 2569 580
rect 2519 497 2569 546
rect 2553 463 2569 497
rect 2519 414 2569 463
rect 2553 380 2569 414
rect 2519 364 2569 380
rect 2217 310 2417 326
rect 2217 276 2371 310
rect 2405 276 2417 310
rect 2217 260 2417 276
rect 1545 177 1887 202
rect 1545 168 1837 177
rect 1821 143 1837 168
rect 1871 143 1887 177
rect 2069 176 2087 210
rect 1266 56 1511 90
rect 1620 118 1769 134
rect 1821 127 1887 143
rect 1933 152 1999 168
rect 1620 84 1636 118
rect 1670 84 1719 118
rect 1753 84 1769 118
rect 1620 17 1769 84
rect 1933 118 1949 152
rect 1983 118 1999 152
rect 1933 17 1999 118
rect 2035 120 2087 176
rect 2069 86 2087 120
rect 2035 70 2087 86
rect 2121 210 2171 226
rect 2155 176 2171 210
rect 2121 120 2171 176
rect 2155 86 2171 120
rect 2121 17 2171 86
rect 2217 190 2283 260
rect 2451 226 2485 364
rect 2417 210 2485 226
rect 2217 156 2233 190
rect 2267 156 2283 190
rect 2217 120 2283 156
rect 2217 86 2233 120
rect 2267 86 2283 120
rect 2217 70 2283 86
rect 2317 190 2383 206
rect 2317 156 2333 190
rect 2367 156 2383 190
rect 2317 120 2383 156
rect 2317 86 2333 120
rect 2367 86 2383 120
rect 2317 17 2383 86
rect 2417 176 2433 210
rect 2467 176 2485 210
rect 2417 120 2485 176
rect 2417 86 2433 120
rect 2467 86 2485 120
rect 2417 70 2485 86
rect 2519 210 2569 226
rect 2553 176 2569 210
rect 2519 120 2569 176
rect 2553 86 2569 120
rect 2519 17 2569 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 1087 316 1121 350
rect 1663 316 1697 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1121 319 1663 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfsbp_2
flabel comment s 872 285 872 285 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 699 308 699 308 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 1663 316 1697 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew
flabel corelocali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2592 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2889368
string GDS_START 2870040
<< end >>
