magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1104 561
rect 28 291 78 527
rect 112 391 162 493
rect 196 425 350 527
rect 636 425 702 527
rect 468 391 518 425
rect 820 391 870 425
rect 112 357 870 391
rect 112 289 170 357
rect 17 215 87 255
rect 121 173 170 289
rect 204 289 652 323
rect 204 215 407 289
rect 441 215 552 255
rect 586 215 652 289
rect 686 289 963 323
rect 997 291 1038 527
rect 686 215 752 289
rect 929 255 963 289
rect 796 215 895 255
rect 929 215 1087 255
rect 104 129 170 173
rect 744 17 778 111
rect 912 17 946 111
rect 0 -17 1104 17
<< obsli1 >>
rect 384 459 602 493
rect 384 425 434 459
rect 552 425 602 459
rect 736 459 954 493
rect 736 425 786 459
rect 904 357 954 459
rect 20 95 70 179
rect 204 129 610 181
rect 644 147 1046 181
rect 204 95 254 129
rect 644 95 710 147
rect 812 145 1046 147
rect 20 51 254 95
rect 292 51 710 95
rect 812 51 878 145
rect 980 51 1046 145
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 929 255 963 289 6 A1
port 1 nsew signal input
rlabel locali s 929 215 1087 255 6 A1
port 1 nsew signal input
rlabel locali s 686 289 963 323 6 A1
port 1 nsew signal input
rlabel locali s 686 215 752 289 6 A1
port 1 nsew signal input
rlabel locali s 796 215 895 255 6 A2
port 2 nsew signal input
rlabel locali s 586 215 652 289 6 B1
port 3 nsew signal input
rlabel locali s 204 289 652 323 6 B1
port 3 nsew signal input
rlabel locali s 204 215 407 289 6 B1
port 3 nsew signal input
rlabel locali s 441 215 552 255 6 B2
port 4 nsew signal input
rlabel locali s 17 215 87 255 6 C1
port 5 nsew signal input
rlabel locali s 820 391 870 425 6 Y
port 6 nsew signal output
rlabel locali s 468 391 518 425 6 Y
port 6 nsew signal output
rlabel locali s 121 173 170 289 6 Y
port 6 nsew signal output
rlabel locali s 112 391 162 493 6 Y
port 6 nsew signal output
rlabel locali s 112 357 870 391 6 Y
port 6 nsew signal output
rlabel locali s 112 289 170 357 6 Y
port 6 nsew signal output
rlabel locali s 104 129 170 173 6 Y
port 6 nsew signal output
rlabel locali s 912 17 946 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 744 17 778 111 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 1104 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 997 291 1038 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 636 425 702 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 196 425 350 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 28 291 78 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1104 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1453250
string GDS_START 1444584
<< end >>
