magic
tech sky130A
magscale 1 2
timestamp 1599588201
<< nwell >>
rect -38 285 2338 582
rect -38 261 394 285
rect 881 261 2338 285
<< pwell >>
rect 43 -2 47 3
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 351 66 381 150
rect 539 119 569 203
rect 611 119 641 203
rect 717 66 817 150
rect 859 66 895 150
rect 1057 47 1087 119
rect 1157 47 1187 119
rect 1263 47 1293 131
rect 1335 47 1365 131
rect 1467 47 1497 175
rect 1562 47 1592 119
rect 1671 47 1701 119
rect 1767 47 1797 131
rect 1916 47 1946 131
rect 1995 47 2025 131
rect 2188 47 2218 177
<< pmoshvt >>
rect 79 297 109 497
rect 166 297 196 497
rect 424 389 454 497
rect 508 389 538 497
rect 590 389 620 497
rect 750 389 780 497
rect 836 389 866 497
rect 1049 413 1079 497
rect 1161 413 1191 497
rect 1245 413 1275 497
rect 1359 413 1389 497
rect 1547 329 1577 497
rect 1642 413 1672 497
rect 1728 413 1758 497
rect 1810 413 1840 497
rect 1916 413 1946 497
rect 2000 413 2030 497
rect 2188 297 2218 497
<< ndiff >>
rect 27 119 79 177
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 177
rect 487 165 539 203
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 129 351 150
rect 299 95 307 129
rect 341 95 351 129
rect 299 66 351 95
rect 381 112 433 150
rect 487 131 495 165
rect 529 131 539 165
rect 487 119 539 131
rect 569 119 611 203
rect 641 195 702 203
rect 641 161 651 195
rect 685 161 702 195
rect 641 150 702 161
rect 641 119 717 150
rect 381 78 391 112
rect 425 78 433 112
rect 381 66 433 78
rect 656 66 717 119
rect 817 66 859 150
rect 895 108 951 150
rect 1417 131 1467 175
rect 1213 119 1263 131
rect 895 74 905 108
rect 939 74 951 108
rect 895 66 951 74
rect 1005 101 1057 119
rect 1005 67 1013 101
rect 1047 67 1057 101
rect 1005 47 1057 67
rect 1087 95 1157 119
rect 1087 61 1113 95
rect 1147 61 1157 95
rect 1087 47 1157 61
rect 1187 47 1263 119
rect 1293 47 1335 131
rect 1365 93 1467 131
rect 1365 59 1399 93
rect 1433 59 1467 93
rect 1365 47 1467 59
rect 1497 119 1547 175
rect 1716 119 1767 131
rect 1497 89 1562 119
rect 1497 55 1507 89
rect 1541 55 1562 89
rect 1497 47 1562 55
rect 1592 93 1671 119
rect 1592 59 1617 93
rect 1651 59 1671 93
rect 1592 47 1671 59
rect 1701 47 1767 119
rect 1797 89 1916 131
rect 1797 55 1817 89
rect 1851 55 1916 89
rect 1797 47 1916 55
rect 1946 47 1995 131
rect 2025 93 2081 131
rect 2025 59 2035 93
rect 2069 59 2081 93
rect 2025 47 2081 59
rect 2136 93 2188 177
rect 2136 59 2144 93
rect 2178 59 2188 93
rect 2136 47 2188 59
rect 2218 143 2270 177
rect 2218 109 2228 143
rect 2262 109 2270 143
rect 2218 47 2270 109
<< pdiff >>
rect 1290 505 1340 517
rect 1290 497 1298 505
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 461 166 497
rect 109 427 122 461
rect 156 427 166 461
rect 109 297 166 427
rect 196 477 249 497
rect 196 443 207 477
rect 241 443 249 477
rect 196 409 249 443
rect 196 375 207 409
rect 241 375 249 409
rect 354 461 424 497
rect 354 427 380 461
rect 414 427 424 461
rect 354 389 424 427
rect 454 462 508 497
rect 454 428 464 462
rect 498 428 508 462
rect 454 389 508 428
rect 538 389 590 497
rect 620 477 750 497
rect 620 443 692 477
rect 726 443 750 477
rect 620 389 750 443
rect 780 389 836 497
rect 866 489 922 497
rect 866 455 876 489
rect 910 455 922 489
rect 866 389 922 455
rect 976 471 1049 497
rect 976 437 1005 471
rect 1039 437 1049 471
rect 976 413 1049 437
rect 1079 483 1161 497
rect 1079 449 1117 483
rect 1151 449 1161 483
rect 1079 413 1161 449
rect 1191 459 1245 497
rect 1191 425 1201 459
rect 1235 425 1245 459
rect 1191 413 1245 425
rect 1275 471 1298 497
rect 1332 497 1340 505
rect 1332 471 1359 497
rect 1275 413 1359 471
rect 1389 459 1441 497
rect 1389 425 1399 459
rect 1433 425 1441 459
rect 1389 413 1441 425
rect 1495 485 1547 497
rect 1495 451 1503 485
rect 1537 451 1547 485
rect 196 297 249 375
rect 1495 329 1547 451
rect 1577 477 1642 497
rect 1577 443 1594 477
rect 1628 443 1642 477
rect 1577 413 1642 443
rect 1672 484 1728 497
rect 1672 450 1684 484
rect 1718 450 1728 484
rect 1672 413 1728 450
rect 1758 413 1810 497
rect 1840 489 1916 497
rect 1840 455 1872 489
rect 1906 455 1916 489
rect 1840 413 1916 455
rect 1946 459 2000 497
rect 1946 425 1956 459
rect 1990 425 2000 459
rect 1946 413 2000 425
rect 2030 485 2082 497
rect 2030 451 2040 485
rect 2074 451 2082 485
rect 2030 413 2082 451
rect 2136 485 2188 497
rect 2136 451 2144 485
rect 2178 451 2188 485
rect 2136 417 2188 451
rect 1577 329 1627 413
rect 2136 383 2144 417
rect 2178 383 2188 417
rect 2136 349 2188 383
rect 2136 315 2144 349
rect 2178 315 2188 349
rect 2136 297 2188 315
rect 2218 449 2270 497
rect 2218 415 2228 449
rect 2262 415 2270 449
rect 2218 381 2270 415
rect 2218 347 2228 381
rect 2262 347 2270 381
rect 2218 297 2270 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 95 341 129
rect 495 131 529 165
rect 651 161 685 195
rect 391 78 425 112
rect 905 74 939 108
rect 1013 67 1047 101
rect 1113 61 1147 95
rect 1399 59 1433 93
rect 1507 55 1541 89
rect 1617 59 1651 93
rect 1817 55 1851 89
rect 2035 59 2069 93
rect 2144 59 2178 93
rect 2228 109 2262 143
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 122 427 156 461
rect 207 443 241 477
rect 207 375 241 409
rect 380 427 414 461
rect 464 428 498 462
rect 692 443 726 477
rect 876 455 910 489
rect 1005 437 1039 471
rect 1117 449 1151 483
rect 1201 425 1235 459
rect 1298 471 1332 505
rect 1399 425 1433 459
rect 1503 451 1537 485
rect 1594 443 1628 477
rect 1684 450 1718 484
rect 1872 455 1906 489
rect 1956 425 1990 459
rect 2040 451 2074 485
rect 2144 451 2178 485
rect 2144 383 2178 417
rect 2144 315 2178 349
rect 2228 415 2262 449
rect 2228 347 2262 381
<< poly >>
rect 79 497 109 523
rect 166 497 196 523
rect 424 497 454 523
rect 508 497 538 523
rect 590 497 620 523
rect 750 497 780 523
rect 836 497 866 523
rect 1049 497 1079 523
rect 1161 497 1191 523
rect 1245 497 1275 523
rect 1359 497 1389 523
rect 1547 497 1577 523
rect 1642 497 1672 523
rect 1728 497 1758 523
rect 1810 497 1840 523
rect 1916 497 1946 523
rect 2000 497 2030 523
rect 2188 497 2218 523
rect 424 357 454 389
rect 508 357 538 389
rect 590 357 620 389
rect 307 327 538 357
rect 580 341 641 357
rect 79 269 109 297
rect 46 265 109 269
rect 166 265 196 297
rect 307 295 381 327
rect 280 279 381 295
rect 580 307 590 341
rect 624 307 641 341
rect 750 337 780 389
rect 836 340 866 389
rect 1049 375 1079 413
rect 1033 365 1099 375
rect 730 336 780 337
rect 728 335 780 336
rect 580 291 641 307
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 280 245 312 279
rect 346 245 381 279
rect 280 229 381 245
rect 151 199 205 215
rect 46 196 109 199
rect 79 177 109 196
rect 163 177 193 199
rect 351 150 381 229
rect 444 275 510 285
rect 444 241 460 275
rect 494 248 510 275
rect 494 241 569 248
rect 444 218 569 241
rect 539 203 569 218
rect 611 203 641 291
rect 726 321 780 335
rect 726 287 736 321
rect 770 287 780 321
rect 726 268 780 287
rect 835 324 895 340
rect 835 290 845 324
rect 879 290 895 324
rect 1033 331 1049 365
rect 1083 331 1099 365
rect 1033 321 1099 331
rect 835 274 895 290
rect 1161 279 1191 413
rect 1245 371 1275 413
rect 1245 353 1317 371
rect 1245 319 1273 353
rect 1307 319 1317 353
rect 1245 303 1317 319
rect 717 150 817 176
rect 859 150 895 274
rect 966 263 1191 279
rect 966 229 981 263
rect 1015 249 1191 263
rect 1015 229 1029 249
rect 966 213 1029 229
rect 999 164 1029 213
rect 1133 191 1187 207
rect 539 93 569 119
rect 611 93 641 119
rect 999 134 1087 164
rect 1133 157 1143 191
rect 1177 157 1187 191
rect 1133 141 1187 157
rect 1057 119 1087 134
rect 1157 119 1187 141
rect 1263 131 1293 303
rect 1359 225 1389 413
rect 1547 314 1577 329
rect 1467 284 1577 314
rect 1467 267 1497 284
rect 1335 209 1389 225
rect 1335 175 1345 209
rect 1379 175 1389 209
rect 1431 251 1497 267
rect 1431 217 1441 251
rect 1475 217 1497 251
rect 1642 279 1672 413
rect 1728 381 1758 413
rect 1714 365 1768 381
rect 1714 331 1724 365
rect 1758 331 1768 365
rect 1714 315 1768 331
rect 1642 267 1688 279
rect 1642 255 1701 267
rect 1642 249 1725 255
rect 1659 239 1725 249
rect 1659 237 1681 239
rect 1431 201 1497 217
rect 1467 175 1497 201
rect 1562 191 1629 207
rect 1335 151 1389 175
rect 1335 131 1365 151
rect 351 51 381 66
rect 717 51 817 66
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 817 51
rect 859 40 895 66
rect 1562 157 1585 191
rect 1619 157 1629 191
rect 1562 141 1629 157
rect 1671 205 1681 237
rect 1715 205 1725 239
rect 1671 189 1725 205
rect 1810 229 1840 413
rect 1916 398 1946 413
rect 1882 387 1946 398
rect 1882 384 1944 387
rect 1882 383 1943 384
rect 1882 381 1942 383
rect 1882 380 1941 381
rect 1882 378 1940 380
rect 1882 377 1939 378
rect 1882 376 1938 377
rect 1882 375 1937 376
rect 1882 374 1936 375
rect 1882 373 1934 374
rect 1882 372 1933 373
rect 1882 371 1931 372
rect 1882 370 1930 371
rect 1882 369 1927 370
rect 1882 368 1924 369
rect 1882 287 1912 368
rect 2000 365 2030 413
rect 1985 364 2037 365
rect 1983 363 2037 364
rect 1981 349 2037 363
rect 1981 315 1991 349
rect 2025 315 2037 349
rect 1981 301 2037 315
rect 1983 300 2037 301
rect 1985 299 2037 300
rect 1882 284 1920 287
rect 1882 283 1923 284
rect 1882 282 1926 283
rect 1882 281 1927 282
rect 1882 280 1929 281
rect 1882 279 1930 280
rect 1882 278 1932 279
rect 1882 277 1933 278
rect 1882 276 1934 277
rect 1882 275 1935 276
rect 1882 273 1936 275
rect 1882 272 1937 273
rect 1882 270 1938 272
rect 1882 269 1939 270
rect 1882 268 1940 269
rect 1885 266 1940 268
rect 1887 265 1941 266
rect 1889 264 1941 265
rect 1891 263 1941 264
rect 1893 262 1961 263
rect 1894 261 1963 262
rect 1895 260 1965 261
rect 1897 259 1965 260
rect 1898 258 1965 259
rect 1899 257 1965 258
rect 1900 256 1965 257
rect 1901 255 1965 256
rect 1902 253 1965 255
rect 1903 252 1965 253
rect 1904 251 1965 252
rect 1905 249 1965 251
rect 1906 247 1965 249
rect 1907 245 1921 247
rect 1908 243 1921 245
rect 1909 240 1921 243
rect 1910 237 1921 240
rect 1810 228 1865 229
rect 1810 227 1867 228
rect 1810 213 1869 227
rect 1810 193 1825 213
rect 1562 119 1592 141
rect 1671 119 1701 189
rect 1767 179 1825 193
rect 1859 179 1869 213
rect 1911 213 1921 237
rect 1955 213 1965 247
rect 1911 197 1965 213
rect 1767 163 1869 179
rect 1767 131 1797 163
rect 1916 131 1946 197
rect 2007 170 2037 299
rect 2188 265 2218 297
rect 2160 249 2218 265
rect 2160 215 2170 249
rect 2204 215 2218 249
rect 2160 199 2218 215
rect 2188 177 2218 199
rect 2005 169 2037 170
rect 2004 168 2037 169
rect 2003 167 2037 168
rect 1995 146 2037 167
rect 1995 131 2025 146
rect 1057 21 1087 47
rect 1157 21 1187 47
rect 1263 21 1293 47
rect 1335 21 1365 47
rect 1467 21 1497 47
rect 1562 21 1592 47
rect 1671 21 1701 47
rect 1767 21 1797 47
rect 1916 21 1946 47
rect 1995 21 2025 47
rect 2188 21 2218 47
<< polycont >>
rect 590 307 624 341
rect 31 215 65 249
rect 161 215 195 249
rect 312 245 346 279
rect 460 241 494 275
rect 736 287 770 321
rect 845 290 879 324
rect 1049 331 1083 365
rect 1273 319 1307 353
rect 981 229 1015 263
rect 1143 157 1177 191
rect 1345 175 1379 209
rect 1441 217 1475 251
rect 1724 331 1758 365
rect 1585 157 1619 191
rect 1681 205 1715 239
rect 1991 315 2025 349
rect 1825 179 1859 213
rect 1921 213 1955 247
rect 2170 215 2204 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 106 461 172 527
rect 106 427 122 461
rect 156 427 172 461
rect 207 477 241 493
rect 18 375 35 409
rect 207 409 241 443
rect 69 375 173 393
rect 18 359 173 375
rect 28 249 98 325
rect 28 215 31 249
rect 65 215 98 249
rect 28 195 98 215
rect 132 265 173 359
rect 293 397 346 493
rect 380 461 430 480
rect 414 427 430 461
rect 380 411 430 427
rect 241 357 263 380
rect 207 346 263 357
rect 132 255 195 265
rect 132 215 161 255
rect 132 199 195 215
rect 132 161 167 199
rect 19 127 167 161
rect 229 135 263 346
rect 297 279 346 397
rect 297 245 312 279
rect 396 291 430 411
rect 464 462 498 527
rect 464 408 498 428
rect 573 357 624 493
rect 692 477 726 493
rect 860 489 926 527
rect 1282 505 1348 527
rect 860 455 876 489
rect 910 455 926 489
rect 981 471 1055 487
rect 692 421 726 443
rect 981 437 1005 471
rect 1039 437 1055 471
rect 1094 483 1167 493
rect 1094 449 1117 483
rect 1151 449 1167 483
rect 981 421 1015 437
rect 1094 427 1167 449
rect 547 341 624 357
rect 547 307 590 341
rect 396 275 494 291
rect 396 252 460 275
rect 297 214 346 245
rect 411 241 460 252
rect 547 271 624 307
rect 658 387 1015 421
rect 411 237 494 241
rect 658 237 692 387
rect 411 199 617 237
rect 411 180 445 199
rect 19 119 69 127
rect 19 85 35 119
rect 203 119 263 135
rect 19 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 263 119
rect 203 69 263 85
rect 307 146 445 180
rect 307 129 341 146
rect 479 131 495 165
rect 529 131 545 165
rect 307 79 341 95
rect 375 78 391 112
rect 425 78 441 112
rect 103 17 169 59
rect 375 17 441 78
rect 479 17 545 131
rect 583 85 617 199
rect 651 203 692 237
rect 736 321 770 337
rect 651 195 685 203
rect 651 135 685 161
rect 736 85 770 287
rect 583 51 770 85
rect 804 324 879 340
rect 804 290 845 324
rect 804 142 879 290
rect 913 179 947 387
rect 1049 365 1065 391
rect 1083 331 1099 357
rect 1049 315 1099 331
rect 981 263 1015 279
rect 981 213 1015 221
rect 1065 207 1099 315
rect 1133 277 1167 427
rect 1201 459 1235 475
rect 1282 471 1298 505
rect 1332 471 1348 505
rect 1475 485 1549 527
rect 1201 421 1235 425
rect 1399 459 1433 475
rect 1475 451 1503 485
rect 1537 451 1549 485
rect 1475 435 1549 451
rect 1594 477 1628 493
rect 1399 421 1433 425
rect 1201 387 1433 421
rect 1594 401 1628 443
rect 1664 484 1838 493
rect 1664 450 1684 484
rect 1718 450 1838 484
rect 1664 425 1838 450
rect 1872 489 1922 527
rect 1906 455 1922 489
rect 2024 485 2090 527
rect 1872 439 1922 455
rect 1956 459 1990 475
rect 1803 423 1838 425
rect 2024 451 2040 485
rect 2074 451 2090 485
rect 2144 485 2194 527
rect 2178 451 2194 485
rect 1803 407 1842 423
rect 1491 367 1628 401
rect 1491 353 1543 367
rect 1257 319 1273 353
rect 1307 319 1543 353
rect 1662 357 1689 391
rect 1723 387 1768 391
rect 1723 365 1774 387
rect 1723 357 1724 365
rect 1662 333 1724 357
rect 1133 251 1475 277
rect 1133 243 1441 251
rect 1065 191 1195 207
rect 913 143 1029 179
rect 804 57 855 142
rect 889 74 905 108
rect 939 74 955 108
rect 889 17 955 74
rect 995 101 1029 143
rect 1065 157 1143 191
rect 1177 157 1195 191
rect 1065 141 1195 157
rect 995 67 1013 101
rect 1047 67 1063 101
rect 1233 95 1267 243
rect 1301 187 1345 209
rect 1379 187 1407 209
rect 1441 201 1475 217
rect 1335 175 1345 187
rect 1335 153 1373 175
rect 1509 167 1543 319
rect 1097 61 1113 95
rect 1147 61 1267 95
rect 1383 93 1449 109
rect 1383 59 1399 93
rect 1433 59 1449 93
rect 1383 17 1449 59
rect 1491 89 1543 167
rect 1577 331 1724 333
rect 1758 331 1774 365
rect 1808 349 1842 407
rect 1956 417 1990 425
rect 2144 417 2194 451
rect 1956 383 2109 417
rect 1577 299 1704 331
rect 1808 315 1991 349
rect 2025 315 2041 349
rect 1577 191 1619 299
rect 1808 297 1842 315
rect 1577 157 1585 191
rect 1681 255 1715 265
rect 1681 184 1715 205
rect 1749 263 1842 297
rect 2075 265 2109 383
rect 2178 383 2194 417
rect 2144 349 2194 383
rect 2178 315 2194 349
rect 2144 299 2194 315
rect 2228 449 2280 465
rect 2262 415 2280 449
rect 2228 381 2280 415
rect 2262 347 2280 381
rect 2228 292 2280 347
rect 2230 289 2280 292
rect 1577 141 1619 157
rect 1749 107 1783 263
rect 2075 259 2204 265
rect 1905 247 1938 255
rect 1825 213 1859 229
rect 1905 213 1921 247
rect 1972 221 2023 255
rect 1955 213 2023 221
rect 1825 173 1859 179
rect 1965 187 2023 213
rect 1825 139 1931 173
rect 1601 93 1783 107
rect 1491 55 1507 89
rect 1541 55 1557 89
rect 1601 59 1617 93
rect 1651 59 1783 93
rect 1601 51 1783 59
rect 1817 89 1851 105
rect 1897 93 1931 139
rect 1965 153 1989 187
rect 1965 127 2023 153
rect 2069 249 2204 259
rect 2069 215 2170 249
rect 2069 199 2204 215
rect 1897 59 2035 93
rect 2069 59 2103 199
rect 2238 159 2280 289
rect 2228 143 2280 159
rect 2262 109 2280 143
rect 2144 93 2178 109
rect 1817 17 1851 55
rect 2144 17 2178 59
rect 2228 53 2280 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 207 375 241 391
rect 207 357 241 375
rect 161 249 195 255
rect 161 221 195 249
rect 1065 365 1099 391
rect 1065 357 1083 365
rect 1083 357 1099 365
rect 981 229 1015 255
rect 981 221 1015 229
rect 1689 357 1723 391
rect 1301 153 1335 187
rect 1373 175 1379 187
rect 1379 175 1407 187
rect 1373 153 1407 175
rect 1681 239 1715 255
rect 1681 221 1715 239
rect 1938 247 1972 255
rect 1938 221 1955 247
rect 1955 221 1972 247
rect 1989 153 2023 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 0 496 2300 527
rect 194 391 254 397
rect 194 357 207 391
rect 241 388 254 391
rect 1053 391 1111 397
rect 1053 388 1065 391
rect 241 360 1065 388
rect 241 357 254 360
rect 194 351 254 357
rect 1053 357 1065 360
rect 1099 388 1111 391
rect 1677 391 1735 397
rect 1677 388 1689 391
rect 1099 360 1689 388
rect 1099 357 1111 360
rect 1053 351 1111 357
rect 1677 357 1689 360
rect 1723 357 1735 391
rect 1677 351 1735 357
rect 149 255 207 261
rect 149 221 161 255
rect 195 252 207 255
rect 969 255 1027 261
rect 969 252 981 255
rect 195 224 981 252
rect 195 221 207 224
rect 149 215 207 221
rect 969 221 981 224
rect 1015 252 1027 255
rect 1669 255 1727 261
rect 1669 252 1681 255
rect 1015 224 1681 252
rect 1015 221 1027 224
rect 969 215 1027 221
rect 1669 221 1681 224
rect 1715 221 1727 255
rect 1669 215 1727 221
rect 1926 255 1984 261
rect 1926 221 1938 255
rect 1972 221 1984 255
rect 1926 193 1984 221
rect 1289 187 1419 193
rect 1289 153 1301 187
rect 1335 153 1373 187
rect 1407 184 1419 187
rect 1926 187 2035 193
rect 1926 184 1989 187
rect 1407 156 1989 184
rect 1407 153 1419 156
rect 1289 147 1419 153
rect 1977 153 1989 156
rect 2023 153 2035 187
rect 1977 147 2035 153
rect 0 17 2300 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
rect 0 -48 2300 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfrtp_1
flabel nwell s 34 528 63 556 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 43 -2 47 3 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel metal1 s 31 534 63 554 0 FreeSans 200 0 0 0 VPWR
port 9 nsew
flabel metal1 s 39 -10 57 7 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel corelocali s 312 289 346 323 0 FreeSans 200 0 0 0 SCE
port 5 nsew
flabel corelocali s 815 289 849 323 0 FreeSans 200 0 0 0 SCD
port 4 nsew
flabel corelocali s 559 289 593 323 0 FreeSans 200 0 0 0 D
port 2 nsew
flabel corelocali s 1965 221 1999 255 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 40 221 74 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 40 289 74 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew
flabel corelocali s 1989 153 2023 187 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew
flabel corelocali s 2234 85 2268 119 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 2234 289 2268 323 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 2234 357 2268 391 0 FreeSans 400 0 0 0 Q
port 10 nsew
flabel corelocali s 2234 425 2268 459 0 FreeSans 400 0 0 0 Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2300 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 157964
string GDS_START 139136
string path 0.000 0.000 11.500 0.000 
<< end >>
