magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 213 356 279 547
rect 21 287 87 356
rect 121 310 279 356
rect 121 184 172 310
rect 409 236 551 356
rect 601 270 670 356
rect 586 184 636 226
rect 121 150 636 184
rect 121 70 172 150
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 123 581 369 615
rect 123 390 179 581
rect 313 492 369 581
rect 409 526 461 649
rect 495 492 561 596
rect 601 526 635 649
rect 675 492 741 596
rect 313 458 741 492
rect 313 390 738 424
rect 20 17 86 226
rect 313 252 355 390
rect 272 218 355 252
rect 704 226 738 390
rect 672 116 738 226
rect 400 17 466 116
rect 500 66 738 116
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel locali s 601 270 670 356 6 A1
port 1 nsew signal input
rlabel locali s 409 236 551 356 6 A2
port 2 nsew signal input
rlabel locali s 21 287 87 356 6 B1
port 3 nsew signal input
rlabel locali s 586 184 636 226 6 Y
port 4 nsew signal output
rlabel locali s 213 356 279 547 6 Y
port 4 nsew signal output
rlabel locali s 121 310 279 356 6 Y
port 4 nsew signal output
rlabel locali s 121 184 172 310 6 Y
port 4 nsew signal output
rlabel locali s 121 150 636 184 6 Y
port 4 nsew signal output
rlabel locali s 121 70 172 150 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 768 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 768 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 4117936
string GDS_START 4111010
<< end >>
