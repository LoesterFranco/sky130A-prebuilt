magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 3718 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 277 47 307 177
rect 361 47 391 177
rect 569 47 599 177
rect 653 47 683 177
rect 757 47 787 177
rect 841 47 871 177
rect 945 47 975 177
rect 1029 47 1059 177
rect 1133 47 1163 177
rect 1217 47 1247 177
rect 1321 47 1351 177
rect 1405 47 1435 177
rect 1613 47 1643 177
rect 1697 47 1727 177
rect 1801 47 1831 177
rect 1885 47 1915 177
rect 2093 47 2123 177
rect 2177 47 2207 177
rect 2281 47 2311 177
rect 2365 47 2395 177
rect 2469 47 2499 177
rect 2553 47 2583 177
rect 2657 47 2687 177
rect 2741 47 2771 177
rect 2845 47 2875 177
rect 2929 47 2959 177
rect 3033 47 3063 177
rect 3117 47 3147 177
rect 3221 47 3251 177
rect 3305 47 3335 177
rect 3409 47 3439 177
rect 3493 47 3523 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 561 297 597 497
rect 655 297 691 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
rect 1605 297 1641 497
rect 1699 297 1735 497
rect 1793 297 1829 497
rect 1887 297 1923 497
rect 2085 297 2121 497
rect 2179 297 2215 497
rect 2273 297 2309 497
rect 2367 297 2403 497
rect 2461 297 2497 497
rect 2555 297 2591 497
rect 2649 297 2685 497
rect 2743 297 2779 497
rect 2837 297 2873 497
rect 2931 297 2967 497
rect 3025 297 3061 497
rect 3119 297 3155 497
rect 3213 297 3249 497
rect 3307 297 3343 497
rect 3401 297 3437 497
rect 3495 297 3531 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 169 173 177
rect 119 135 129 169
rect 163 135 173 169
rect 119 47 173 135
rect 203 93 277 177
rect 203 59 223 93
rect 257 59 277 93
rect 203 47 277 59
rect 307 169 361 177
rect 307 135 317 169
rect 351 135 361 169
rect 307 47 361 135
rect 391 94 453 177
rect 391 60 411 94
rect 445 60 453 94
rect 391 47 453 60
rect 507 94 569 177
rect 507 60 515 94
rect 549 60 569 94
rect 507 47 569 60
rect 599 169 653 177
rect 599 135 609 169
rect 643 135 653 169
rect 599 101 653 135
rect 599 67 609 101
rect 643 67 653 101
rect 599 47 653 67
rect 683 93 757 177
rect 683 59 703 93
rect 737 59 757 93
rect 683 47 757 59
rect 787 169 841 177
rect 787 135 797 169
rect 831 135 841 169
rect 787 101 841 135
rect 787 67 797 101
rect 831 67 841 101
rect 787 47 841 67
rect 871 165 945 177
rect 871 131 891 165
rect 925 131 945 165
rect 871 93 945 131
rect 871 59 891 93
rect 925 59 945 93
rect 871 47 945 59
rect 975 169 1029 177
rect 975 135 985 169
rect 1019 135 1029 169
rect 975 101 1029 135
rect 975 67 985 101
rect 1019 67 1029 101
rect 975 47 1029 67
rect 1059 165 1133 177
rect 1059 131 1079 165
rect 1113 131 1133 165
rect 1059 93 1133 131
rect 1059 59 1079 93
rect 1113 59 1133 93
rect 1059 47 1133 59
rect 1163 169 1217 177
rect 1163 135 1173 169
rect 1207 135 1217 169
rect 1163 101 1217 135
rect 1163 67 1173 101
rect 1207 67 1217 101
rect 1163 47 1217 67
rect 1247 93 1321 177
rect 1247 59 1267 93
rect 1301 59 1321 93
rect 1247 47 1321 59
rect 1351 169 1405 177
rect 1351 135 1361 169
rect 1395 135 1405 169
rect 1351 101 1405 135
rect 1351 67 1361 101
rect 1395 67 1405 101
rect 1351 47 1405 67
rect 1435 94 1497 177
rect 1435 60 1455 94
rect 1489 60 1497 94
rect 1435 47 1497 60
rect 1551 94 1613 177
rect 1551 60 1559 94
rect 1593 60 1613 94
rect 1551 47 1613 60
rect 1643 169 1697 177
rect 1643 135 1653 169
rect 1687 135 1697 169
rect 1643 47 1697 135
rect 1727 93 1801 177
rect 1727 59 1747 93
rect 1781 59 1801 93
rect 1727 47 1801 59
rect 1831 169 1885 177
rect 1831 135 1841 169
rect 1875 135 1885 169
rect 1831 47 1885 135
rect 1915 165 1977 177
rect 1915 131 1935 165
rect 1969 131 1977 165
rect 1915 97 1977 131
rect 1915 63 1935 97
rect 1969 63 1977 97
rect 1915 47 1977 63
rect 2031 165 2093 177
rect 2031 131 2039 165
rect 2073 131 2093 165
rect 2031 93 2093 131
rect 2031 59 2039 93
rect 2073 59 2093 93
rect 2031 47 2093 59
rect 2123 169 2177 177
rect 2123 135 2133 169
rect 2167 135 2177 169
rect 2123 101 2177 135
rect 2123 67 2133 101
rect 2167 67 2177 101
rect 2123 47 2177 67
rect 2207 93 2281 177
rect 2207 59 2227 93
rect 2261 59 2281 93
rect 2207 47 2281 59
rect 2311 169 2365 177
rect 2311 135 2321 169
rect 2355 135 2365 169
rect 2311 101 2365 135
rect 2311 67 2321 101
rect 2355 67 2365 101
rect 2311 47 2365 67
rect 2395 93 2469 177
rect 2395 59 2415 93
rect 2449 59 2469 93
rect 2395 47 2469 59
rect 2499 169 2553 177
rect 2499 135 2509 169
rect 2543 135 2553 169
rect 2499 101 2553 135
rect 2499 67 2509 101
rect 2543 67 2553 101
rect 2499 47 2553 67
rect 2583 93 2657 177
rect 2583 59 2603 93
rect 2637 59 2657 93
rect 2583 47 2657 59
rect 2687 169 2741 177
rect 2687 135 2697 169
rect 2731 135 2741 169
rect 2687 101 2741 135
rect 2687 67 2697 101
rect 2731 67 2741 101
rect 2687 47 2741 67
rect 2771 94 2845 177
rect 2771 60 2791 94
rect 2825 60 2845 94
rect 2771 47 2845 60
rect 2875 169 2929 177
rect 2875 135 2885 169
rect 2919 135 2929 169
rect 2875 101 2929 135
rect 2875 67 2885 101
rect 2919 67 2929 101
rect 2875 47 2929 67
rect 2959 93 3033 177
rect 2959 59 2979 93
rect 3013 59 3033 93
rect 2959 47 3033 59
rect 3063 169 3117 177
rect 3063 135 3073 169
rect 3107 135 3117 169
rect 3063 101 3117 135
rect 3063 67 3073 101
rect 3107 67 3117 101
rect 3063 47 3117 67
rect 3147 93 3221 177
rect 3147 59 3167 93
rect 3201 59 3221 93
rect 3147 47 3221 59
rect 3251 169 3305 177
rect 3251 135 3261 169
rect 3295 135 3305 169
rect 3251 101 3305 135
rect 3251 67 3261 101
rect 3295 67 3305 101
rect 3251 47 3305 67
rect 3335 93 3409 177
rect 3335 59 3355 93
rect 3389 59 3409 93
rect 3335 47 3409 59
rect 3439 169 3493 177
rect 3439 135 3449 169
rect 3483 135 3493 169
rect 3439 101 3493 135
rect 3439 67 3449 101
rect 3483 67 3493 101
rect 3439 47 3493 67
rect 3523 165 3585 177
rect 3523 131 3543 165
rect 3577 131 3585 165
rect 3523 93 3585 131
rect 3523 59 3543 93
rect 3577 59 3585 93
rect 3523 47 3585 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 417 175 497
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 417 363 497
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 453 497
rect 399 451 411 485
rect 445 451 453 485
rect 399 417 453 451
rect 399 383 411 417
rect 445 383 453 417
rect 399 349 453 383
rect 399 315 411 349
rect 445 315 453 349
rect 399 297 453 315
rect 507 485 561 497
rect 507 451 515 485
rect 549 451 561 485
rect 507 417 561 451
rect 507 383 515 417
rect 549 383 561 417
rect 507 349 561 383
rect 507 315 515 349
rect 549 315 561 349
rect 507 297 561 315
rect 597 485 655 497
rect 597 451 609 485
rect 643 451 655 485
rect 597 417 655 451
rect 597 383 609 417
rect 643 383 655 417
rect 597 349 655 383
rect 597 315 609 349
rect 643 315 655 349
rect 597 297 655 315
rect 691 485 749 497
rect 691 451 703 485
rect 737 451 749 485
rect 691 417 749 451
rect 691 383 703 417
rect 737 383 749 417
rect 691 297 749 383
rect 785 485 843 497
rect 785 451 797 485
rect 831 451 843 485
rect 785 417 843 451
rect 785 383 797 417
rect 831 383 843 417
rect 785 349 843 383
rect 785 315 797 349
rect 831 315 843 349
rect 785 297 843 315
rect 879 485 937 497
rect 879 451 891 485
rect 925 451 937 485
rect 879 417 937 451
rect 879 383 891 417
rect 925 383 937 417
rect 879 349 937 383
rect 879 315 891 349
rect 925 315 937 349
rect 879 297 937 315
rect 973 485 1031 497
rect 973 451 985 485
rect 1019 451 1031 485
rect 973 417 1031 451
rect 973 383 985 417
rect 1019 383 1031 417
rect 973 349 1031 383
rect 973 315 985 349
rect 1019 315 1031 349
rect 973 297 1031 315
rect 1067 485 1125 497
rect 1067 451 1079 485
rect 1113 451 1125 485
rect 1067 417 1125 451
rect 1067 383 1079 417
rect 1113 383 1125 417
rect 1067 349 1125 383
rect 1067 315 1079 349
rect 1113 315 1125 349
rect 1067 297 1125 315
rect 1161 485 1219 497
rect 1161 451 1173 485
rect 1207 451 1219 485
rect 1161 417 1219 451
rect 1161 383 1173 417
rect 1207 383 1219 417
rect 1161 349 1219 383
rect 1161 315 1173 349
rect 1207 315 1219 349
rect 1161 297 1219 315
rect 1255 485 1313 497
rect 1255 451 1267 485
rect 1301 451 1313 485
rect 1255 417 1313 451
rect 1255 383 1267 417
rect 1301 383 1313 417
rect 1255 297 1313 383
rect 1349 485 1407 497
rect 1349 451 1361 485
rect 1395 451 1407 485
rect 1349 417 1407 451
rect 1349 383 1361 417
rect 1395 383 1407 417
rect 1349 349 1407 383
rect 1349 315 1361 349
rect 1395 315 1407 349
rect 1349 297 1407 315
rect 1443 485 1497 497
rect 1443 451 1455 485
rect 1489 451 1497 485
rect 1443 417 1497 451
rect 1443 383 1455 417
rect 1489 383 1497 417
rect 1443 349 1497 383
rect 1443 315 1455 349
rect 1489 315 1497 349
rect 1443 297 1497 315
rect 1551 485 1605 497
rect 1551 451 1559 485
rect 1593 451 1605 485
rect 1551 417 1605 451
rect 1551 383 1559 417
rect 1593 383 1605 417
rect 1551 349 1605 383
rect 1551 315 1559 349
rect 1593 315 1605 349
rect 1551 297 1605 315
rect 1641 417 1699 497
rect 1641 383 1653 417
rect 1687 383 1699 417
rect 1641 349 1699 383
rect 1641 315 1653 349
rect 1687 315 1699 349
rect 1641 297 1699 315
rect 1735 485 1793 497
rect 1735 451 1747 485
rect 1781 451 1793 485
rect 1735 417 1793 451
rect 1735 383 1747 417
rect 1781 383 1793 417
rect 1735 297 1793 383
rect 1829 417 1887 497
rect 1829 383 1841 417
rect 1875 383 1887 417
rect 1829 349 1887 383
rect 1829 315 1841 349
rect 1875 315 1887 349
rect 1829 297 1887 315
rect 1923 485 1977 497
rect 1923 451 1935 485
rect 1969 451 1977 485
rect 1923 417 1977 451
rect 1923 383 1935 417
rect 1969 383 1977 417
rect 1923 349 1977 383
rect 1923 315 1935 349
rect 1969 315 1977 349
rect 1923 297 1977 315
rect 2031 485 2085 497
rect 2031 451 2039 485
rect 2073 451 2085 485
rect 2031 417 2085 451
rect 2031 383 2039 417
rect 2073 383 2085 417
rect 2031 349 2085 383
rect 2031 315 2039 349
rect 2073 315 2085 349
rect 2031 297 2085 315
rect 2121 485 2179 497
rect 2121 451 2133 485
rect 2167 451 2179 485
rect 2121 417 2179 451
rect 2121 383 2133 417
rect 2167 383 2179 417
rect 2121 349 2179 383
rect 2121 315 2133 349
rect 2167 315 2179 349
rect 2121 297 2179 315
rect 2215 485 2273 497
rect 2215 451 2227 485
rect 2261 451 2273 485
rect 2215 417 2273 451
rect 2215 383 2227 417
rect 2261 383 2273 417
rect 2215 297 2273 383
rect 2309 485 2367 497
rect 2309 451 2321 485
rect 2355 451 2367 485
rect 2309 417 2367 451
rect 2309 383 2321 417
rect 2355 383 2367 417
rect 2309 349 2367 383
rect 2309 315 2321 349
rect 2355 315 2367 349
rect 2309 297 2367 315
rect 2403 485 2461 497
rect 2403 451 2415 485
rect 2449 451 2461 485
rect 2403 417 2461 451
rect 2403 383 2415 417
rect 2449 383 2461 417
rect 2403 297 2461 383
rect 2497 485 2555 497
rect 2497 451 2509 485
rect 2543 451 2555 485
rect 2497 417 2555 451
rect 2497 383 2509 417
rect 2543 383 2555 417
rect 2497 349 2555 383
rect 2497 315 2509 349
rect 2543 315 2555 349
rect 2497 297 2555 315
rect 2591 485 2649 497
rect 2591 451 2603 485
rect 2637 451 2649 485
rect 2591 417 2649 451
rect 2591 383 2603 417
rect 2637 383 2649 417
rect 2591 297 2649 383
rect 2685 485 2743 497
rect 2685 451 2697 485
rect 2731 451 2743 485
rect 2685 417 2743 451
rect 2685 383 2697 417
rect 2731 383 2743 417
rect 2685 349 2743 383
rect 2685 315 2697 349
rect 2731 315 2743 349
rect 2685 297 2743 315
rect 2779 485 2837 497
rect 2779 451 2791 485
rect 2825 451 2837 485
rect 2779 417 2837 451
rect 2779 383 2791 417
rect 2825 383 2837 417
rect 2779 297 2837 383
rect 2873 485 2931 497
rect 2873 451 2885 485
rect 2919 451 2931 485
rect 2873 417 2931 451
rect 2873 383 2885 417
rect 2919 383 2931 417
rect 2873 349 2931 383
rect 2873 315 2885 349
rect 2919 315 2931 349
rect 2873 297 2931 315
rect 2967 485 3025 497
rect 2967 451 2979 485
rect 3013 451 3025 485
rect 2967 417 3025 451
rect 2967 383 2979 417
rect 3013 383 3025 417
rect 2967 297 3025 383
rect 3061 485 3119 497
rect 3061 451 3073 485
rect 3107 451 3119 485
rect 3061 417 3119 451
rect 3061 383 3073 417
rect 3107 383 3119 417
rect 3061 349 3119 383
rect 3061 315 3073 349
rect 3107 315 3119 349
rect 3061 297 3119 315
rect 3155 485 3213 497
rect 3155 451 3167 485
rect 3201 451 3213 485
rect 3155 417 3213 451
rect 3155 383 3167 417
rect 3201 383 3213 417
rect 3155 297 3213 383
rect 3249 485 3307 497
rect 3249 451 3261 485
rect 3295 451 3307 485
rect 3249 417 3307 451
rect 3249 383 3261 417
rect 3295 383 3307 417
rect 3249 349 3307 383
rect 3249 315 3261 349
rect 3295 315 3307 349
rect 3249 297 3307 315
rect 3343 485 3401 497
rect 3343 451 3355 485
rect 3389 451 3401 485
rect 3343 417 3401 451
rect 3343 383 3355 417
rect 3389 383 3401 417
rect 3343 297 3401 383
rect 3437 485 3495 497
rect 3437 451 3449 485
rect 3483 451 3495 485
rect 3437 417 3495 451
rect 3437 383 3449 417
rect 3483 383 3495 417
rect 3437 349 3495 383
rect 3437 315 3449 349
rect 3483 315 3495 349
rect 3437 297 3495 315
rect 3531 485 3585 497
rect 3531 451 3543 485
rect 3577 451 3585 485
rect 3531 417 3585 451
rect 3531 383 3543 417
rect 3577 383 3585 417
rect 3531 349 3585 383
rect 3531 315 3543 349
rect 3577 315 3585 349
rect 3531 297 3585 315
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 135 163 169
rect 223 59 257 93
rect 317 135 351 169
rect 411 60 445 94
rect 515 60 549 94
rect 609 135 643 169
rect 609 67 643 101
rect 703 59 737 93
rect 797 135 831 169
rect 797 67 831 101
rect 891 131 925 165
rect 891 59 925 93
rect 985 135 1019 169
rect 985 67 1019 101
rect 1079 131 1113 165
rect 1079 59 1113 93
rect 1173 135 1207 169
rect 1173 67 1207 101
rect 1267 59 1301 93
rect 1361 135 1395 169
rect 1361 67 1395 101
rect 1455 60 1489 94
rect 1559 60 1593 94
rect 1653 135 1687 169
rect 1747 59 1781 93
rect 1841 135 1875 169
rect 1935 131 1969 165
rect 1935 63 1969 97
rect 2039 131 2073 165
rect 2039 59 2073 93
rect 2133 135 2167 169
rect 2133 67 2167 101
rect 2227 59 2261 93
rect 2321 135 2355 169
rect 2321 67 2355 101
rect 2415 59 2449 93
rect 2509 135 2543 169
rect 2509 67 2543 101
rect 2603 59 2637 93
rect 2697 135 2731 169
rect 2697 67 2731 101
rect 2791 60 2825 94
rect 2885 135 2919 169
rect 2885 67 2919 101
rect 2979 59 3013 93
rect 3073 135 3107 169
rect 3073 67 3107 101
rect 3167 59 3201 93
rect 3261 135 3295 169
rect 3261 67 3295 101
rect 3355 59 3389 93
rect 3449 135 3483 169
rect 3449 67 3483 101
rect 3543 131 3577 165
rect 3543 59 3577 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 411 315 445 349
rect 515 451 549 485
rect 515 383 549 417
rect 515 315 549 349
rect 609 451 643 485
rect 609 383 643 417
rect 609 315 643 349
rect 703 451 737 485
rect 703 383 737 417
rect 797 451 831 485
rect 797 383 831 417
rect 797 315 831 349
rect 891 451 925 485
rect 891 383 925 417
rect 891 315 925 349
rect 985 451 1019 485
rect 985 383 1019 417
rect 985 315 1019 349
rect 1079 451 1113 485
rect 1079 383 1113 417
rect 1079 315 1113 349
rect 1173 451 1207 485
rect 1173 383 1207 417
rect 1173 315 1207 349
rect 1267 451 1301 485
rect 1267 383 1301 417
rect 1361 451 1395 485
rect 1361 383 1395 417
rect 1361 315 1395 349
rect 1455 451 1489 485
rect 1455 383 1489 417
rect 1455 315 1489 349
rect 1559 451 1593 485
rect 1559 383 1593 417
rect 1559 315 1593 349
rect 1653 383 1687 417
rect 1653 315 1687 349
rect 1747 451 1781 485
rect 1747 383 1781 417
rect 1841 383 1875 417
rect 1841 315 1875 349
rect 1935 451 1969 485
rect 1935 383 1969 417
rect 1935 315 1969 349
rect 2039 451 2073 485
rect 2039 383 2073 417
rect 2039 315 2073 349
rect 2133 451 2167 485
rect 2133 383 2167 417
rect 2133 315 2167 349
rect 2227 451 2261 485
rect 2227 383 2261 417
rect 2321 451 2355 485
rect 2321 383 2355 417
rect 2321 315 2355 349
rect 2415 451 2449 485
rect 2415 383 2449 417
rect 2509 451 2543 485
rect 2509 383 2543 417
rect 2509 315 2543 349
rect 2603 451 2637 485
rect 2603 383 2637 417
rect 2697 451 2731 485
rect 2697 383 2731 417
rect 2697 315 2731 349
rect 2791 451 2825 485
rect 2791 383 2825 417
rect 2885 451 2919 485
rect 2885 383 2919 417
rect 2885 315 2919 349
rect 2979 451 3013 485
rect 2979 383 3013 417
rect 3073 451 3107 485
rect 3073 383 3107 417
rect 3073 315 3107 349
rect 3167 451 3201 485
rect 3167 383 3201 417
rect 3261 451 3295 485
rect 3261 383 3295 417
rect 3261 315 3295 349
rect 3355 451 3389 485
rect 3355 383 3389 417
rect 3449 451 3483 485
rect 3449 383 3483 417
rect 3449 315 3483 349
rect 3543 451 3577 485
rect 3543 383 3577 417
rect 3543 315 3577 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 561 497 597 523
rect 655 497 691 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 1605 497 1641 523
rect 1699 497 1735 523
rect 1793 497 1829 523
rect 1887 497 1923 523
rect 2085 497 2121 523
rect 2179 497 2215 523
rect 2273 497 2309 523
rect 2367 497 2403 523
rect 2461 497 2497 523
rect 2555 497 2591 523
rect 2649 497 2685 523
rect 2743 497 2779 523
rect 2837 497 2873 523
rect 2931 497 2967 523
rect 3025 497 3061 523
rect 3119 497 3155 523
rect 3213 497 3249 523
rect 3307 497 3343 523
rect 3401 497 3437 523
rect 3495 497 3531 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 561 282 597 297
rect 655 282 691 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 1605 282 1641 297
rect 1699 282 1735 297
rect 1793 282 1829 297
rect 1887 282 1923 297
rect 2085 282 2121 297
rect 2179 282 2215 297
rect 2273 282 2309 297
rect 2367 282 2403 297
rect 2461 282 2497 297
rect 2555 282 2591 297
rect 2649 282 2685 297
rect 2743 282 2779 297
rect 2837 282 2873 297
rect 2931 282 2967 297
rect 3025 282 3061 297
rect 3119 282 3155 297
rect 3213 282 3249 297
rect 3307 282 3343 297
rect 3401 282 3437 297
rect 3495 282 3531 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 79 249 401 265
rect 79 215 129 249
rect 163 215 197 249
rect 231 215 265 249
rect 299 215 333 249
rect 367 215 401 249
rect 79 199 401 215
rect 559 265 599 282
rect 653 265 693 282
rect 747 265 787 282
rect 841 265 881 282
rect 935 265 975 282
rect 1029 265 1069 282
rect 559 249 1069 265
rect 559 215 601 249
rect 635 215 669 249
rect 703 215 737 249
rect 771 215 805 249
rect 839 215 1069 249
rect 559 199 1069 215
rect 1123 265 1163 282
rect 1217 265 1257 282
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 1123 249 1445 265
rect 1123 215 1165 249
rect 1199 215 1233 249
rect 1267 215 1301 249
rect 1335 215 1369 249
rect 1403 215 1445 249
rect 1123 199 1445 215
rect 1603 265 1643 282
rect 1697 265 1737 282
rect 1791 265 1831 282
rect 1885 265 1925 282
rect 1603 249 1925 265
rect 1603 215 1637 249
rect 1671 215 1705 249
rect 1739 215 1773 249
rect 1807 215 1841 249
rect 1875 215 1925 249
rect 1603 199 1925 215
rect 2083 265 2123 282
rect 2177 265 2217 282
rect 2271 265 2311 282
rect 2365 265 2405 282
rect 2459 265 2499 282
rect 2553 265 2593 282
rect 2647 265 2687 282
rect 2741 265 2781 282
rect 2835 265 2875 282
rect 2929 265 2969 282
rect 3023 265 3063 282
rect 3117 265 3157 282
rect 3211 265 3251 282
rect 3305 265 3345 282
rect 3399 265 3439 282
rect 3493 265 3533 282
rect 2083 249 3533 265
rect 2083 215 2099 249
rect 2133 215 2167 249
rect 2201 215 2235 249
rect 2269 215 2303 249
rect 2337 215 2371 249
rect 2405 215 2439 249
rect 2473 215 2507 249
rect 2541 215 2575 249
rect 2609 215 2643 249
rect 2677 215 2711 249
rect 2745 215 2779 249
rect 2813 215 2847 249
rect 2881 215 2915 249
rect 2949 215 2983 249
rect 3017 215 3051 249
rect 3085 215 3119 249
rect 3153 215 3187 249
rect 3221 215 3255 249
rect 3289 215 3323 249
rect 3357 215 3533 249
rect 2083 199 3533 215
rect 89 177 119 199
rect 173 177 203 199
rect 277 177 307 199
rect 361 177 391 199
rect 569 177 599 199
rect 653 177 683 199
rect 757 177 787 199
rect 841 177 871 199
rect 945 177 975 199
rect 1029 177 1059 199
rect 1133 177 1163 199
rect 1217 177 1247 199
rect 1321 177 1351 199
rect 1405 177 1435 199
rect 1613 177 1643 199
rect 1697 177 1727 199
rect 1801 177 1831 199
rect 1885 177 1915 199
rect 2093 177 2123 199
rect 2177 177 2207 199
rect 2281 177 2311 199
rect 2365 177 2395 199
rect 2469 177 2499 199
rect 2553 177 2583 199
rect 2657 177 2687 199
rect 2741 177 2771 199
rect 2845 177 2875 199
rect 2929 177 2959 199
rect 3033 177 3063 199
rect 3117 177 3147 199
rect 3221 177 3251 199
rect 3305 177 3335 199
rect 3409 177 3439 199
rect 3493 177 3523 199
rect 89 21 119 47
rect 173 21 203 47
rect 277 21 307 47
rect 361 21 391 47
rect 569 21 599 47
rect 653 21 683 47
rect 757 21 787 47
rect 841 21 871 47
rect 945 21 975 47
rect 1029 21 1059 47
rect 1133 21 1163 47
rect 1217 21 1247 47
rect 1321 21 1351 47
rect 1405 21 1435 47
rect 1613 21 1643 47
rect 1697 21 1727 47
rect 1801 21 1831 47
rect 1885 21 1915 47
rect 2093 21 2123 47
rect 2177 21 2207 47
rect 2281 21 2311 47
rect 2365 21 2395 47
rect 2469 21 2499 47
rect 2553 21 2583 47
rect 2657 21 2687 47
rect 2741 21 2771 47
rect 2845 21 2875 47
rect 2929 21 2959 47
rect 3033 21 3063 47
rect 3117 21 3147 47
rect 3221 21 3251 47
rect 3305 21 3335 47
rect 3409 21 3439 47
rect 3493 21 3523 47
<< polycont >>
rect 129 215 163 249
rect 197 215 231 249
rect 265 215 299 249
rect 333 215 367 249
rect 601 215 635 249
rect 669 215 703 249
rect 737 215 771 249
rect 805 215 839 249
rect 1165 215 1199 249
rect 1233 215 1267 249
rect 1301 215 1335 249
rect 1369 215 1403 249
rect 1637 215 1671 249
rect 1705 215 1739 249
rect 1773 215 1807 249
rect 1841 215 1875 249
rect 2099 215 2133 249
rect 2167 215 2201 249
rect 2235 215 2269 249
rect 2303 215 2337 249
rect 2371 215 2405 249
rect 2439 215 2473 249
rect 2507 215 2541 249
rect 2575 215 2609 249
rect 2643 215 2677 249
rect 2711 215 2745 249
rect 2779 215 2813 249
rect 2847 215 2881 249
rect 2915 215 2949 249
rect 2983 215 3017 249
rect 3051 215 3085 249
rect 3119 215 3153 249
rect 3187 215 3221 249
rect 3255 215 3289 249
rect 3323 215 3357 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 19 485 461 493
rect 19 451 35 485
rect 69 459 223 485
rect 69 451 79 459
rect 19 417 79 451
rect 213 451 223 459
rect 257 459 411 485
rect 257 451 267 459
rect 19 383 35 417
rect 69 383 79 417
rect 19 349 79 383
rect 19 315 35 349
rect 69 315 79 349
rect 19 165 79 315
rect 113 417 179 425
rect 113 357 129 417
rect 163 357 179 417
rect 213 417 267 451
rect 401 451 411 459
rect 445 451 461 485
rect 213 383 223 417
rect 257 383 267 417
rect 213 367 267 383
rect 301 417 367 425
rect 113 349 179 357
rect 113 315 129 349
rect 163 333 179 349
rect 301 357 317 417
rect 351 357 367 417
rect 301 349 367 357
rect 301 333 317 349
rect 163 315 317 333
rect 351 315 367 349
rect 113 299 367 315
rect 401 417 461 451
rect 401 383 411 417
rect 445 383 461 417
rect 401 349 461 383
rect 401 315 411 349
rect 445 315 461 349
rect 401 299 461 315
rect 505 485 559 527
rect 505 451 515 485
rect 549 451 559 485
rect 505 417 559 451
rect 505 383 515 417
rect 549 383 559 417
rect 505 349 559 383
rect 505 315 515 349
rect 549 315 559 349
rect 505 299 559 315
rect 593 485 659 493
rect 593 425 609 485
rect 643 425 659 485
rect 593 417 659 425
rect 593 383 609 417
rect 643 383 659 417
rect 593 349 659 383
rect 693 485 747 527
rect 693 451 703 485
rect 737 451 747 485
rect 693 417 747 451
rect 693 383 703 417
rect 737 383 747 417
rect 693 367 747 383
rect 781 485 847 493
rect 781 425 797 485
rect 831 425 847 485
rect 781 417 847 425
rect 781 383 797 417
rect 831 383 847 417
rect 593 315 609 349
rect 643 333 659 349
rect 781 349 847 383
rect 781 333 797 349
rect 643 315 797 333
rect 831 315 847 349
rect 593 299 847 315
rect 881 485 935 527
rect 881 451 891 485
rect 925 451 935 485
rect 881 417 935 451
rect 881 383 891 417
rect 925 383 935 417
rect 881 349 935 383
rect 881 315 891 349
rect 925 315 935 349
rect 881 299 935 315
rect 969 485 1035 493
rect 969 451 985 485
rect 1019 451 1035 485
rect 969 417 1035 451
rect 969 383 985 417
rect 1019 383 1035 417
rect 969 349 1035 383
rect 969 315 985 349
rect 1019 315 1035 349
rect 969 265 1035 315
rect 1069 485 1123 527
rect 1069 451 1079 485
rect 1113 451 1123 485
rect 1069 417 1123 451
rect 1069 383 1079 417
rect 1113 383 1123 417
rect 1069 349 1123 383
rect 1069 315 1079 349
rect 1113 315 1123 349
rect 1069 299 1123 315
rect 1157 485 1223 493
rect 1157 451 1173 485
rect 1207 451 1223 485
rect 1157 417 1223 451
rect 1157 357 1173 417
rect 1207 357 1223 417
rect 1257 485 1311 527
rect 1257 451 1267 485
rect 1301 451 1311 485
rect 1257 417 1311 451
rect 1257 383 1267 417
rect 1301 383 1311 417
rect 1257 367 1311 383
rect 1345 485 1411 493
rect 1345 451 1361 485
rect 1395 451 1411 485
rect 1345 417 1411 451
rect 1157 349 1223 357
rect 1157 315 1173 349
rect 1207 333 1223 349
rect 1345 357 1361 417
rect 1395 357 1411 417
rect 1345 349 1411 357
rect 1345 333 1361 349
rect 1207 315 1361 333
rect 1395 315 1411 349
rect 1157 299 1411 315
rect 1445 485 1499 527
rect 1445 451 1455 485
rect 1489 451 1499 485
rect 1445 417 1499 451
rect 1445 383 1455 417
rect 1489 383 1499 417
rect 1445 349 1499 383
rect 1445 315 1455 349
rect 1489 315 1499 349
rect 1445 299 1499 315
rect 1543 485 1985 493
rect 1543 451 1559 485
rect 1593 459 1747 485
rect 1593 451 1603 459
rect 1543 417 1603 451
rect 1737 451 1747 459
rect 1781 459 1935 485
rect 1781 451 1791 459
rect 1543 383 1559 417
rect 1593 383 1603 417
rect 1543 349 1603 383
rect 1543 315 1559 349
rect 1593 315 1603 349
rect 1543 299 1603 315
rect 1637 417 1703 425
rect 1637 357 1653 417
rect 1687 357 1703 417
rect 1737 417 1791 451
rect 1925 451 1935 459
rect 1969 451 1985 485
rect 1737 383 1747 417
rect 1781 383 1791 417
rect 1737 367 1791 383
rect 1825 417 1891 425
rect 1637 349 1703 357
rect 1637 315 1653 349
rect 1687 333 1703 349
rect 1825 357 1841 417
rect 1875 357 1891 417
rect 1825 349 1891 357
rect 1825 333 1841 349
rect 1687 315 1841 333
rect 1875 315 1891 349
rect 1637 299 1891 315
rect 1925 417 1985 451
rect 1925 383 1935 417
rect 1969 383 1985 417
rect 1925 349 1985 383
rect 1925 315 1935 349
rect 1969 315 1985 349
rect 1925 265 1985 315
rect 2029 485 2083 527
rect 2029 451 2039 485
rect 2073 451 2083 485
rect 2029 417 2083 451
rect 2029 383 2039 417
rect 2073 383 2083 417
rect 2029 349 2083 383
rect 2029 315 2039 349
rect 2073 315 2083 349
rect 2029 299 2083 315
rect 2117 485 2183 493
rect 2117 451 2133 485
rect 2167 451 2183 485
rect 2117 417 2183 451
rect 2117 383 2133 417
rect 2167 383 2183 417
rect 2117 349 2183 383
rect 2217 485 2271 527
rect 2217 451 2227 485
rect 2261 451 2271 485
rect 2217 417 2271 451
rect 2217 383 2227 417
rect 2261 383 2271 417
rect 2217 367 2271 383
rect 2305 485 2371 493
rect 2305 451 2321 485
rect 2355 451 2371 485
rect 2305 417 2371 451
rect 2305 383 2321 417
rect 2355 383 2371 417
rect 2117 315 2133 349
rect 2167 333 2183 349
rect 2305 349 2371 383
rect 2405 485 2459 527
rect 2405 451 2415 485
rect 2449 451 2459 485
rect 2405 417 2459 451
rect 2405 383 2415 417
rect 2449 383 2459 417
rect 2405 367 2459 383
rect 2493 485 2559 493
rect 2493 451 2509 485
rect 2543 451 2559 485
rect 2493 417 2559 451
rect 2493 383 2509 417
rect 2543 383 2559 417
rect 2305 333 2321 349
rect 2167 315 2321 333
rect 2355 333 2371 349
rect 2493 349 2559 383
rect 2593 485 2647 527
rect 2593 451 2603 485
rect 2637 451 2647 485
rect 2593 417 2647 451
rect 2593 383 2603 417
rect 2637 383 2647 417
rect 2593 367 2647 383
rect 2681 485 2747 493
rect 2681 451 2697 485
rect 2731 451 2747 485
rect 2681 417 2747 451
rect 2681 383 2697 417
rect 2731 383 2747 417
rect 2493 333 2509 349
rect 2355 315 2509 333
rect 2543 333 2559 349
rect 2681 349 2747 383
rect 2781 485 2835 527
rect 2781 451 2791 485
rect 2825 451 2835 485
rect 2781 417 2835 451
rect 2781 383 2791 417
rect 2825 383 2835 417
rect 2781 367 2835 383
rect 2869 485 2935 493
rect 2869 451 2885 485
rect 2919 451 2935 485
rect 2869 417 2935 451
rect 2869 383 2885 417
rect 2919 383 2935 417
rect 2681 333 2697 349
rect 2543 315 2697 333
rect 2731 333 2747 349
rect 2869 349 2935 383
rect 2969 485 3023 527
rect 2969 451 2979 485
rect 3013 451 3023 485
rect 2969 417 3023 451
rect 2969 383 2979 417
rect 3013 383 3023 417
rect 2969 367 3023 383
rect 3057 485 3123 493
rect 3057 451 3073 485
rect 3107 451 3123 485
rect 3057 417 3123 451
rect 3057 383 3073 417
rect 3107 383 3123 417
rect 2869 333 2885 349
rect 2731 315 2885 333
rect 2919 333 2935 349
rect 3057 349 3123 383
rect 3157 485 3211 527
rect 3157 451 3167 485
rect 3201 451 3211 485
rect 3157 417 3211 451
rect 3157 383 3167 417
rect 3201 383 3211 417
rect 3157 367 3211 383
rect 3245 485 3311 493
rect 3245 451 3261 485
rect 3295 451 3311 485
rect 3245 417 3311 451
rect 3245 383 3261 417
rect 3295 383 3311 417
rect 3057 333 3073 349
rect 2919 315 3073 333
rect 3107 333 3123 349
rect 3245 349 3311 383
rect 3345 485 3399 527
rect 3345 451 3355 485
rect 3389 451 3399 485
rect 3345 417 3399 451
rect 3345 383 3355 417
rect 3389 383 3399 417
rect 3345 367 3399 383
rect 3433 485 3499 493
rect 3433 451 3449 485
rect 3483 451 3499 485
rect 3433 417 3499 451
rect 3433 383 3449 417
rect 3483 383 3499 417
rect 3245 333 3261 349
rect 3107 315 3261 333
rect 3295 333 3311 349
rect 3433 349 3499 383
rect 3433 333 3449 349
rect 3295 315 3449 333
rect 3483 315 3499 349
rect 2117 299 3499 315
rect 3533 485 3587 527
rect 3533 451 3543 485
rect 3577 451 3587 485
rect 3533 417 3587 451
rect 3533 383 3543 417
rect 3577 383 3587 417
rect 3533 349 3587 383
rect 3533 315 3543 349
rect 3577 315 3587 349
rect 3533 299 3587 315
rect 113 249 383 265
rect 113 215 129 249
rect 163 215 197 249
rect 231 215 265 249
rect 299 215 333 249
rect 367 215 383 249
rect 585 249 855 265
rect 585 215 601 249
rect 635 215 669 249
rect 703 215 737 249
rect 771 215 805 249
rect 839 215 855 249
rect 969 249 1419 265
rect 969 215 1165 249
rect 1199 215 1233 249
rect 1267 215 1301 249
rect 1335 215 1369 249
rect 1403 215 1419 249
rect 1621 249 1891 265
rect 1621 215 1637 249
rect 1671 215 1705 249
rect 1739 215 1773 249
rect 1807 215 1841 249
rect 1875 215 1891 249
rect 1925 249 3373 265
rect 1925 215 2099 249
rect 2133 215 2167 249
rect 2201 215 2235 249
rect 2269 215 2303 249
rect 2337 215 2371 249
rect 2405 215 2439 249
rect 2473 215 2507 249
rect 2541 215 2575 249
rect 2609 215 2643 249
rect 2677 215 2711 249
rect 2745 215 2779 249
rect 2813 215 2847 249
rect 2881 215 2915 249
rect 2949 215 2983 249
rect 3017 215 3051 249
rect 3085 215 3119 249
rect 3153 215 3187 249
rect 3221 215 3255 249
rect 3289 215 3323 249
rect 3357 215 3373 249
rect 19 131 35 165
rect 69 131 79 165
rect 19 119 79 131
rect 113 169 847 181
rect 113 135 129 169
rect 163 145 317 169
rect 163 135 179 145
rect 113 119 179 135
rect 301 135 317 145
rect 351 145 609 169
rect 351 135 367 145
rect 301 119 367 135
rect 593 135 609 145
rect 643 145 797 169
rect 643 135 659 145
rect 19 63 35 119
rect 69 85 79 119
rect 213 93 267 109
rect 213 85 223 93
rect 69 63 223 85
rect 19 59 223 63
rect 257 85 267 93
rect 401 94 461 110
rect 401 85 411 94
rect 257 60 411 85
rect 445 60 461 94
rect 257 59 461 60
rect 19 51 461 59
rect 505 94 559 110
rect 505 60 515 94
rect 549 60 559 94
rect 505 17 559 60
rect 593 101 659 135
rect 781 135 797 145
rect 831 135 847 169
rect 593 67 609 101
rect 643 67 659 101
rect 593 51 659 67
rect 693 93 747 109
rect 693 59 703 93
rect 737 59 747 93
rect 693 17 747 59
rect 781 101 847 135
rect 781 67 797 101
rect 831 67 847 101
rect 781 51 847 67
rect 881 165 935 181
rect 881 131 891 165
rect 925 131 935 165
rect 881 93 935 131
rect 881 59 891 93
rect 925 59 935 93
rect 881 17 935 59
rect 969 169 1035 215
rect 969 135 985 169
rect 1019 135 1035 169
rect 969 101 1035 135
rect 969 67 985 101
rect 1019 67 1035 101
rect 969 51 1035 67
rect 1069 165 1123 181
rect 1069 131 1079 165
rect 1113 131 1123 165
rect 1069 93 1123 131
rect 1069 59 1079 93
rect 1113 59 1123 93
rect 1069 17 1123 59
rect 1157 169 1891 181
rect 1157 135 1173 169
rect 1207 145 1361 169
rect 1207 135 1223 145
rect 1157 101 1223 135
rect 1345 135 1361 145
rect 1395 145 1653 169
rect 1395 135 1411 145
rect 1157 67 1173 101
rect 1207 67 1223 101
rect 1157 51 1223 67
rect 1257 93 1311 109
rect 1257 59 1267 93
rect 1301 59 1311 93
rect 1257 17 1311 59
rect 1345 101 1411 135
rect 1637 135 1653 145
rect 1687 145 1841 169
rect 1687 135 1703 145
rect 1637 119 1703 135
rect 1825 135 1841 145
rect 1875 135 1891 169
rect 1825 119 1891 135
rect 1925 165 1985 215
rect 3417 181 3499 299
rect 1925 131 1935 165
rect 1969 131 1985 165
rect 1925 119 1985 131
rect 1345 67 1361 101
rect 1395 67 1411 101
rect 1345 51 1411 67
rect 1445 94 1499 110
rect 1445 60 1455 94
rect 1489 60 1499 94
rect 1445 17 1499 60
rect 1543 94 1603 110
rect 1543 60 1559 94
rect 1593 85 1603 94
rect 1737 93 1791 109
rect 1737 85 1747 93
rect 1593 60 1747 85
rect 1543 59 1747 60
rect 1781 85 1791 93
rect 1925 85 1935 119
rect 1781 63 1935 85
rect 1969 63 1985 119
rect 1781 59 1985 63
rect 1543 51 1985 59
rect 2029 165 2083 181
rect 2029 131 2039 165
rect 2073 131 2083 165
rect 2029 93 2083 131
rect 2029 59 2039 93
rect 2073 59 2083 93
rect 2029 17 2083 59
rect 2117 169 3499 181
rect 2117 135 2133 169
rect 2167 145 2321 169
rect 2167 135 2183 145
rect 2117 101 2183 135
rect 2305 135 2321 145
rect 2355 145 2509 169
rect 2355 135 2371 145
rect 2117 67 2133 101
rect 2167 67 2183 101
rect 2117 51 2183 67
rect 2217 93 2271 109
rect 2217 59 2227 93
rect 2261 59 2271 93
rect 2217 17 2271 59
rect 2305 101 2371 135
rect 2493 135 2509 145
rect 2543 145 2697 169
rect 2543 135 2559 145
rect 2305 67 2321 101
rect 2355 67 2371 101
rect 2305 51 2371 67
rect 2405 93 2459 109
rect 2405 59 2415 93
rect 2449 59 2459 93
rect 2405 17 2459 59
rect 2493 101 2559 135
rect 2681 135 2697 145
rect 2731 145 2885 169
rect 2731 135 2747 145
rect 2493 67 2509 101
rect 2543 67 2559 101
rect 2493 51 2559 67
rect 2593 93 2647 109
rect 2593 59 2603 93
rect 2637 59 2647 93
rect 2593 17 2647 59
rect 2681 101 2747 135
rect 2869 135 2885 145
rect 2919 145 3073 169
rect 2919 135 2935 145
rect 2681 67 2697 101
rect 2731 67 2747 101
rect 2681 51 2747 67
rect 2781 94 2835 110
rect 2781 60 2791 94
rect 2825 60 2835 94
rect 2781 17 2835 60
rect 2869 101 2935 135
rect 3057 135 3073 145
rect 3107 145 3261 169
rect 3107 135 3123 145
rect 2869 67 2885 101
rect 2919 67 2935 101
rect 2869 51 2935 67
rect 2969 93 3023 109
rect 2969 59 2979 93
rect 3013 59 3023 93
rect 2969 17 3023 59
rect 3057 101 3123 135
rect 3245 135 3261 145
rect 3295 145 3449 169
rect 3295 135 3311 145
rect 3057 67 3073 101
rect 3107 67 3123 101
rect 3057 51 3123 67
rect 3157 93 3211 109
rect 3157 59 3167 93
rect 3201 59 3211 93
rect 3157 17 3211 59
rect 3245 101 3311 135
rect 3433 135 3449 145
rect 3483 135 3499 169
rect 3245 67 3261 101
rect 3295 67 3311 101
rect 3245 51 3311 67
rect 3345 93 3399 109
rect 3345 59 3355 93
rect 3389 59 3399 93
rect 3345 17 3399 59
rect 3433 101 3499 135
rect 3433 67 3449 101
rect 3483 67 3499 101
rect 3433 51 3499 67
rect 3533 165 3587 181
rect 3533 131 3543 165
rect 3577 131 3587 165
rect 3533 93 3587 131
rect 3533 59 3543 93
rect 3577 59 3587 93
rect 3533 17 3587 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 3341 527 3375 561
rect 3433 527 3467 561
rect 3525 527 3559 561
rect 3617 527 3651 561
rect 129 383 163 391
rect 129 357 163 383
rect 317 383 351 391
rect 317 357 351 383
rect 609 451 643 459
rect 609 425 643 451
rect 797 451 831 459
rect 797 425 831 451
rect 1173 383 1207 391
rect 1173 357 1207 383
rect 1361 383 1395 391
rect 1361 357 1395 383
rect 1653 383 1687 391
rect 1653 357 1687 383
rect 1841 383 1875 391
rect 1841 357 1875 383
rect 35 97 69 119
rect 35 85 69 97
rect 1935 97 1969 119
rect 1935 85 1969 97
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
rect 3341 -17 3375 17
rect 3433 -17 3467 17
rect 3525 -17 3559 17
rect 3617 -17 3651 17
<< metal1 >>
rect 0 561 3680 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3680 561
rect 0 496 3680 527
rect 597 459 655 465
rect 597 425 609 459
rect 643 456 655 459
rect 785 459 843 465
rect 785 456 797 459
rect 643 428 797 456
rect 643 425 655 428
rect 597 419 655 425
rect 785 425 797 428
rect 831 456 843 459
rect 831 428 1532 456
rect 831 425 843 428
rect 785 419 843 425
rect 117 391 175 397
rect 117 357 129 391
rect 163 388 175 391
rect 305 391 363 397
rect 305 388 317 391
rect 163 360 317 388
rect 163 357 175 360
rect 117 351 175 357
rect 305 357 317 360
rect 351 388 363 391
rect 1161 391 1219 397
rect 1161 388 1173 391
rect 351 360 1173 388
rect 351 357 363 360
rect 305 351 363 357
rect 1161 357 1173 360
rect 1207 388 1219 391
rect 1349 391 1407 397
rect 1349 388 1361 391
rect 1207 360 1361 388
rect 1207 357 1219 360
rect 1161 351 1219 357
rect 1349 357 1361 360
rect 1395 357 1407 391
rect 1504 388 1532 428
rect 1641 391 1699 397
rect 1641 388 1653 391
rect 1504 360 1653 388
rect 1349 351 1407 357
rect 1641 357 1653 360
rect 1687 388 1699 391
rect 1829 391 1887 397
rect 1829 388 1841 391
rect 1687 360 1841 388
rect 1687 357 1699 360
rect 1641 351 1699 357
rect 1829 357 1841 360
rect 1875 357 1887 391
rect 1829 351 1887 357
rect 23 119 81 125
rect 23 85 35 119
rect 69 116 81 119
rect 1923 119 1981 125
rect 1923 116 1935 119
rect 69 88 1935 116
rect 69 85 81 88
rect 23 79 81 85
rect 1923 85 1935 88
rect 1969 85 1981 119
rect 1923 79 1981 85
rect 0 17 3680 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3680 17
rect 0 -48 3680 -17
<< labels >>
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel corelocali s 3433 221 3467 255 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 703 221 737 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel corelocali s 213 221 247 255 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 1777 221 1811 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
rlabel comment s 0 0 0 0 4 mux2_16
<< properties >>
string FIXED_BBOX 0 0 3680 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3430384
string GDS_START 3403082
<< end >>
