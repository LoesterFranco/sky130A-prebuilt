magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 117 324 503 358
rect 117 233 183 324
rect 231 236 297 290
rect 369 270 503 324
rect 605 404 639 547
rect 605 370 937 404
rect 697 236 829 310
rect 231 202 829 236
rect 871 168 937 370
rect 666 134 937 168
rect 666 119 732 134
rect 871 70 937 134
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 460 89 649
rect 213 426 263 596
rect 309 494 359 596
rect 399 528 465 649
rect 499 581 735 615
rect 499 494 565 581
rect 309 460 565 494
rect 49 392 571 426
rect 49 168 83 392
rect 537 336 571 392
rect 679 472 735 581
rect 769 506 835 649
rect 869 472 937 596
rect 679 438 937 472
rect 537 270 625 336
rect 49 134 244 168
rect 23 17 142 100
rect 178 70 244 134
rect 278 17 344 168
rect 394 134 632 168
rect 394 70 460 134
rect 496 17 564 100
rect 598 85 632 134
rect 768 85 835 100
rect 598 51 835 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel locali s 369 270 503 324 6 A
port 1 nsew signal input
rlabel locali s 117 324 503 358 6 A
port 1 nsew signal input
rlabel locali s 117 233 183 324 6 A
port 1 nsew signal input
rlabel locali s 697 236 829 310 6 B
port 2 nsew signal input
rlabel locali s 231 236 297 290 6 B
port 2 nsew signal input
rlabel locali s 231 202 829 236 6 B
port 2 nsew signal input
rlabel locali s 871 168 937 370 6 X
port 3 nsew signal output
rlabel locali s 871 70 937 134 6 X
port 3 nsew signal output
rlabel locali s 666 134 937 168 6 X
port 3 nsew signal output
rlabel locali s 666 119 732 134 6 X
port 3 nsew signal output
rlabel locali s 605 404 639 547 6 X
port 3 nsew signal output
rlabel locali s 605 370 937 404 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 960 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 558652
string GDS_START 550956
<< end >>
