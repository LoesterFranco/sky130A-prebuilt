magic
tech sky130A
magscale 1 2
timestamp 1599588218
<< nwell >>
rect -38 332 2630 704
<< pwell >>
rect 0 0 2592 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 558 368 594 592
rect 648 368 684 592
rect 738 368 774 592
rect 828 368 864 592
rect 920 368 956 592
rect 1010 368 1046 592
rect 1102 368 1138 592
rect 1192 368 1228 592
rect 1292 368 1328 592
rect 1382 368 1418 592
rect 1472 368 1508 592
rect 1562 368 1598 592
rect 1652 368 1688 592
rect 1742 368 1778 592
rect 1832 368 1868 592
rect 1922 368 1958 592
rect 2012 368 2048 592
rect 2102 368 2138 592
rect 2192 368 2228 592
rect 2282 368 2318 592
rect 2372 368 2408 592
rect 2472 368 2508 592
<< nmoslvt >>
rect 87 74 117 222
rect 173 74 203 222
rect 259 74 289 222
rect 346 74 376 222
rect 558 74 588 222
rect 644 74 674 222
rect 744 74 774 222
rect 830 74 860 222
rect 930 74 960 222
rect 1016 74 1046 222
rect 1102 74 1132 222
rect 1188 74 1218 222
rect 1274 74 1304 222
rect 1360 74 1390 222
rect 1446 74 1476 222
rect 1532 74 1562 222
rect 1632 74 1662 222
rect 1718 74 1748 222
rect 1818 74 1848 222
rect 1904 74 1934 222
rect 2004 74 2034 222
rect 2090 74 2120 222
rect 2190 74 2220 222
rect 2276 74 2306 222
rect 2378 74 2408 222
rect 2464 74 2494 222
<< ndiff >>
rect 30 210 87 222
rect 30 176 42 210
rect 76 176 87 210
rect 30 120 87 176
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 142 173 222
rect 117 108 128 142
rect 162 108 173 142
rect 117 74 173 108
rect 203 210 259 222
rect 203 176 214 210
rect 248 176 259 210
rect 203 120 259 176
rect 203 86 214 120
rect 248 86 259 120
rect 203 74 259 86
rect 289 142 346 222
rect 289 108 300 142
rect 334 108 346 142
rect 289 74 346 108
rect 376 210 433 222
rect 376 176 387 210
rect 421 176 433 210
rect 376 120 433 176
rect 376 86 387 120
rect 421 86 433 120
rect 376 74 433 86
rect 487 210 558 222
rect 487 176 499 210
rect 533 176 558 210
rect 487 120 558 176
rect 487 86 499 120
rect 533 86 558 120
rect 487 74 558 86
rect 588 210 644 222
rect 588 176 599 210
rect 633 176 644 210
rect 588 120 644 176
rect 588 86 599 120
rect 633 86 644 120
rect 588 74 644 86
rect 674 146 744 222
rect 674 112 685 146
rect 719 112 744 146
rect 674 74 744 112
rect 774 210 830 222
rect 774 176 785 210
rect 819 176 830 210
rect 774 120 830 176
rect 774 86 785 120
rect 819 86 830 120
rect 774 74 830 86
rect 860 146 930 222
rect 860 112 871 146
rect 905 112 930 146
rect 860 74 930 112
rect 960 210 1016 222
rect 960 176 971 210
rect 1005 176 1016 210
rect 960 120 1016 176
rect 960 86 971 120
rect 1005 86 1016 120
rect 960 74 1016 86
rect 1046 210 1102 222
rect 1046 176 1057 210
rect 1091 176 1102 210
rect 1046 133 1102 176
rect 1046 99 1057 133
rect 1091 99 1102 133
rect 1046 74 1102 99
rect 1132 210 1188 222
rect 1132 176 1143 210
rect 1177 176 1188 210
rect 1132 120 1188 176
rect 1132 86 1143 120
rect 1177 86 1188 120
rect 1132 74 1188 86
rect 1218 210 1274 222
rect 1218 176 1229 210
rect 1263 176 1274 210
rect 1218 120 1274 176
rect 1218 86 1229 120
rect 1263 86 1274 120
rect 1218 74 1274 86
rect 1304 210 1360 222
rect 1304 176 1315 210
rect 1349 176 1360 210
rect 1304 120 1360 176
rect 1304 86 1315 120
rect 1349 86 1360 120
rect 1304 74 1360 86
rect 1390 210 1446 222
rect 1390 176 1401 210
rect 1435 176 1446 210
rect 1390 120 1446 176
rect 1390 86 1401 120
rect 1435 86 1446 120
rect 1390 74 1446 86
rect 1476 210 1532 222
rect 1476 176 1487 210
rect 1521 176 1532 210
rect 1476 120 1532 176
rect 1476 86 1487 120
rect 1521 86 1532 120
rect 1476 74 1532 86
rect 1562 210 1632 222
rect 1562 176 1573 210
rect 1607 176 1632 210
rect 1562 120 1632 176
rect 1562 86 1573 120
rect 1607 86 1632 120
rect 1562 74 1632 86
rect 1662 210 1718 222
rect 1662 176 1673 210
rect 1707 176 1718 210
rect 1662 120 1718 176
rect 1662 86 1673 120
rect 1707 86 1718 120
rect 1662 74 1718 86
rect 1748 210 1818 222
rect 1748 176 1759 210
rect 1793 176 1818 210
rect 1748 120 1818 176
rect 1748 86 1759 120
rect 1793 86 1818 120
rect 1748 74 1818 86
rect 1848 210 1904 222
rect 1848 176 1859 210
rect 1893 176 1904 210
rect 1848 120 1904 176
rect 1848 86 1859 120
rect 1893 86 1904 120
rect 1848 74 1904 86
rect 1934 210 2004 222
rect 1934 176 1945 210
rect 1979 176 2004 210
rect 1934 120 2004 176
rect 1934 86 1945 120
rect 1979 86 2004 120
rect 1934 74 2004 86
rect 2034 210 2090 222
rect 2034 176 2045 210
rect 2079 176 2090 210
rect 2034 120 2090 176
rect 2034 86 2045 120
rect 2079 86 2090 120
rect 2034 74 2090 86
rect 2120 210 2190 222
rect 2120 176 2131 210
rect 2165 176 2190 210
rect 2120 120 2190 176
rect 2120 86 2131 120
rect 2165 86 2190 120
rect 2120 74 2190 86
rect 2220 210 2276 222
rect 2220 176 2231 210
rect 2265 176 2276 210
rect 2220 120 2276 176
rect 2220 86 2231 120
rect 2265 86 2276 120
rect 2220 74 2276 86
rect 2306 210 2378 222
rect 2306 176 2317 210
rect 2351 176 2378 210
rect 2306 120 2378 176
rect 2306 86 2317 120
rect 2351 86 2378 120
rect 2306 74 2378 86
rect 2408 210 2464 222
rect 2408 176 2419 210
rect 2453 176 2464 210
rect 2408 120 2464 176
rect 2408 86 2419 120
rect 2453 86 2464 120
rect 2408 74 2464 86
rect 2494 210 2565 222
rect 2494 176 2519 210
rect 2553 176 2565 210
rect 2494 120 2565 176
rect 2494 86 2519 120
rect 2553 86 2565 120
rect 2494 74 2565 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 440 83 476
rect 27 406 39 440
rect 73 406 83 440
rect 27 368 83 406
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 508 173 546
rect 119 474 129 508
rect 163 474 173 508
rect 119 368 173 474
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 497 263 546
rect 209 463 219 497
rect 253 463 263 497
rect 209 414 263 463
rect 209 380 219 414
rect 253 380 263 414
rect 209 368 263 380
rect 299 580 353 592
rect 299 546 309 580
rect 343 546 353 580
rect 299 478 353 546
rect 299 444 309 478
rect 343 444 353 478
rect 299 368 353 444
rect 389 580 445 592
rect 389 546 399 580
rect 433 546 445 580
rect 389 497 445 546
rect 389 463 399 497
rect 433 463 445 497
rect 389 414 445 463
rect 389 380 399 414
rect 433 380 445 414
rect 389 368 445 380
rect 502 580 558 592
rect 502 546 514 580
rect 548 546 558 580
rect 502 497 558 546
rect 502 463 514 497
rect 548 463 558 497
rect 502 414 558 463
rect 502 380 514 414
rect 548 380 558 414
rect 502 368 558 380
rect 594 580 648 592
rect 594 546 604 580
rect 638 546 648 580
rect 594 497 648 546
rect 594 463 604 497
rect 638 463 648 497
rect 594 414 648 463
rect 594 380 604 414
rect 638 380 648 414
rect 594 368 648 380
rect 684 580 738 592
rect 684 546 694 580
rect 728 546 738 580
rect 684 482 738 546
rect 684 448 694 482
rect 728 448 738 482
rect 684 368 738 448
rect 774 580 828 592
rect 774 546 784 580
rect 818 546 828 580
rect 774 497 828 546
rect 774 463 784 497
rect 818 463 828 497
rect 774 414 828 463
rect 774 380 784 414
rect 818 380 828 414
rect 774 368 828 380
rect 864 580 920 592
rect 864 546 874 580
rect 908 546 920 580
rect 864 482 920 546
rect 864 448 874 482
rect 908 448 920 482
rect 864 368 920 448
rect 956 580 1010 592
rect 956 546 966 580
rect 1000 546 1010 580
rect 956 497 1010 546
rect 956 463 966 497
rect 1000 463 1010 497
rect 956 414 1010 463
rect 956 380 966 414
rect 1000 380 1010 414
rect 956 368 1010 380
rect 1046 580 1102 592
rect 1046 546 1056 580
rect 1090 546 1102 580
rect 1046 503 1102 546
rect 1046 469 1056 503
rect 1090 469 1102 503
rect 1046 435 1102 469
rect 1046 401 1056 435
rect 1090 401 1102 435
rect 1046 368 1102 401
rect 1138 580 1192 592
rect 1138 546 1148 580
rect 1182 546 1192 580
rect 1138 497 1192 546
rect 1138 463 1148 497
rect 1182 463 1192 497
rect 1138 419 1192 463
rect 1138 385 1148 419
rect 1182 385 1192 419
rect 1138 368 1192 385
rect 1228 580 1292 592
rect 1228 546 1248 580
rect 1282 546 1292 580
rect 1228 482 1292 546
rect 1228 448 1248 482
rect 1282 448 1292 482
rect 1228 368 1292 448
rect 1328 580 1382 592
rect 1328 546 1338 580
rect 1372 546 1382 580
rect 1328 497 1382 546
rect 1328 463 1338 497
rect 1372 463 1382 497
rect 1328 418 1382 463
rect 1328 384 1338 418
rect 1372 384 1382 418
rect 1328 368 1382 384
rect 1418 580 1472 592
rect 1418 546 1428 580
rect 1462 546 1472 580
rect 1418 482 1472 546
rect 1418 448 1428 482
rect 1462 448 1472 482
rect 1418 368 1472 448
rect 1508 580 1562 592
rect 1508 546 1518 580
rect 1552 546 1562 580
rect 1508 497 1562 546
rect 1508 463 1518 497
rect 1552 463 1562 497
rect 1508 418 1562 463
rect 1508 384 1518 418
rect 1552 384 1562 418
rect 1508 368 1562 384
rect 1598 580 1652 592
rect 1598 546 1608 580
rect 1642 546 1652 580
rect 1598 503 1652 546
rect 1598 469 1608 503
rect 1642 469 1652 503
rect 1598 435 1652 469
rect 1598 401 1608 435
rect 1642 401 1652 435
rect 1598 368 1652 401
rect 1688 580 1742 592
rect 1688 546 1698 580
rect 1732 546 1742 580
rect 1688 497 1742 546
rect 1688 463 1698 497
rect 1732 463 1742 497
rect 1688 418 1742 463
rect 1688 384 1698 418
rect 1732 384 1742 418
rect 1688 368 1742 384
rect 1778 580 1832 592
rect 1778 546 1788 580
rect 1822 546 1832 580
rect 1778 503 1832 546
rect 1778 469 1788 503
rect 1822 469 1832 503
rect 1778 435 1832 469
rect 1778 401 1788 435
rect 1822 401 1832 435
rect 1778 368 1832 401
rect 1868 580 1922 592
rect 1868 546 1878 580
rect 1912 546 1922 580
rect 1868 497 1922 546
rect 1868 463 1878 497
rect 1912 463 1922 497
rect 1868 418 1922 463
rect 1868 384 1878 418
rect 1912 384 1922 418
rect 1868 368 1922 384
rect 1958 580 2012 592
rect 1958 546 1968 580
rect 2002 546 2012 580
rect 1958 503 2012 546
rect 1958 469 1968 503
rect 2002 469 2012 503
rect 1958 435 2012 469
rect 1958 401 1968 435
rect 2002 401 2012 435
rect 1958 368 2012 401
rect 2048 580 2102 592
rect 2048 546 2058 580
rect 2092 546 2102 580
rect 2048 497 2102 546
rect 2048 463 2058 497
rect 2092 463 2102 497
rect 2048 418 2102 463
rect 2048 384 2058 418
rect 2092 384 2102 418
rect 2048 368 2102 384
rect 2138 580 2192 592
rect 2138 546 2148 580
rect 2182 546 2192 580
rect 2138 503 2192 546
rect 2138 469 2148 503
rect 2182 469 2192 503
rect 2138 435 2192 469
rect 2138 401 2148 435
rect 2182 401 2192 435
rect 2138 368 2192 401
rect 2228 580 2282 592
rect 2228 546 2238 580
rect 2272 546 2282 580
rect 2228 497 2282 546
rect 2228 463 2238 497
rect 2272 463 2282 497
rect 2228 418 2282 463
rect 2228 384 2238 418
rect 2272 384 2282 418
rect 2228 368 2282 384
rect 2318 580 2372 592
rect 2318 546 2328 580
rect 2362 546 2372 580
rect 2318 503 2372 546
rect 2318 469 2328 503
rect 2362 469 2372 503
rect 2318 435 2372 469
rect 2318 401 2328 435
rect 2362 401 2372 435
rect 2318 368 2372 401
rect 2408 580 2472 592
rect 2408 546 2428 580
rect 2462 546 2472 580
rect 2408 497 2472 546
rect 2408 463 2428 497
rect 2462 463 2472 497
rect 2408 414 2472 463
rect 2408 380 2428 414
rect 2462 380 2472 414
rect 2408 368 2472 380
rect 2508 580 2564 592
rect 2508 546 2518 580
rect 2552 546 2564 580
rect 2508 497 2564 546
rect 2508 463 2518 497
rect 2552 463 2564 497
rect 2508 414 2564 463
rect 2508 380 2518 414
rect 2552 380 2564 414
rect 2508 368 2564 380
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 128 108 162 142
rect 214 176 248 210
rect 214 86 248 120
rect 300 108 334 142
rect 387 176 421 210
rect 387 86 421 120
rect 499 176 533 210
rect 499 86 533 120
rect 599 176 633 210
rect 599 86 633 120
rect 685 112 719 146
rect 785 176 819 210
rect 785 86 819 120
rect 871 112 905 146
rect 971 176 1005 210
rect 971 86 1005 120
rect 1057 176 1091 210
rect 1057 99 1091 133
rect 1143 176 1177 210
rect 1143 86 1177 120
rect 1229 176 1263 210
rect 1229 86 1263 120
rect 1315 176 1349 210
rect 1315 86 1349 120
rect 1401 176 1435 210
rect 1401 86 1435 120
rect 1487 176 1521 210
rect 1487 86 1521 120
rect 1573 176 1607 210
rect 1573 86 1607 120
rect 1673 176 1707 210
rect 1673 86 1707 120
rect 1759 176 1793 210
rect 1759 86 1793 120
rect 1859 176 1893 210
rect 1859 86 1893 120
rect 1945 176 1979 210
rect 1945 86 1979 120
rect 2045 176 2079 210
rect 2045 86 2079 120
rect 2131 176 2165 210
rect 2131 86 2165 120
rect 2231 176 2265 210
rect 2231 86 2265 120
rect 2317 176 2351 210
rect 2317 86 2351 120
rect 2419 176 2453 210
rect 2419 86 2453 120
rect 2519 176 2553 210
rect 2519 86 2553 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 474 163 508
rect 219 546 253 580
rect 219 463 253 497
rect 219 380 253 414
rect 309 546 343 580
rect 309 444 343 478
rect 399 546 433 580
rect 399 463 433 497
rect 399 380 433 414
rect 514 546 548 580
rect 514 463 548 497
rect 514 380 548 414
rect 604 546 638 580
rect 604 463 638 497
rect 604 380 638 414
rect 694 546 728 580
rect 694 448 728 482
rect 784 546 818 580
rect 784 463 818 497
rect 784 380 818 414
rect 874 546 908 580
rect 874 448 908 482
rect 966 546 1000 580
rect 966 463 1000 497
rect 966 380 1000 414
rect 1056 546 1090 580
rect 1056 469 1090 503
rect 1056 401 1090 435
rect 1148 546 1182 580
rect 1148 463 1182 497
rect 1148 385 1182 419
rect 1248 546 1282 580
rect 1248 448 1282 482
rect 1338 546 1372 580
rect 1338 463 1372 497
rect 1338 384 1372 418
rect 1428 546 1462 580
rect 1428 448 1462 482
rect 1518 546 1552 580
rect 1518 463 1552 497
rect 1518 384 1552 418
rect 1608 546 1642 580
rect 1608 469 1642 503
rect 1608 401 1642 435
rect 1698 546 1732 580
rect 1698 463 1732 497
rect 1698 384 1732 418
rect 1788 546 1822 580
rect 1788 469 1822 503
rect 1788 401 1822 435
rect 1878 546 1912 580
rect 1878 463 1912 497
rect 1878 384 1912 418
rect 1968 546 2002 580
rect 1968 469 2002 503
rect 1968 401 2002 435
rect 2058 546 2092 580
rect 2058 463 2092 497
rect 2058 384 2092 418
rect 2148 546 2182 580
rect 2148 469 2182 503
rect 2148 401 2182 435
rect 2238 546 2272 580
rect 2238 463 2272 497
rect 2238 384 2272 418
rect 2328 546 2362 580
rect 2328 469 2362 503
rect 2328 401 2362 435
rect 2428 546 2462 580
rect 2428 463 2462 497
rect 2428 380 2462 414
rect 2518 546 2552 580
rect 2518 463 2552 497
rect 2518 380 2552 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 558 592 594 618
rect 648 592 684 618
rect 738 592 774 618
rect 828 592 864 618
rect 920 592 956 618
rect 1010 592 1046 618
rect 1102 592 1138 618
rect 1192 592 1228 618
rect 1292 592 1328 618
rect 1382 592 1418 618
rect 1472 592 1508 618
rect 1562 592 1598 618
rect 1652 592 1688 618
rect 1742 592 1778 618
rect 1832 592 1868 618
rect 1922 592 1958 618
rect 2012 592 2048 618
rect 2102 592 2138 618
rect 2192 592 2228 618
rect 2282 592 2318 618
rect 2372 592 2408 618
rect 2472 592 2508 618
rect 83 326 119 368
rect 35 310 119 326
rect 35 276 51 310
rect 85 276 119 310
rect 35 260 119 276
rect 173 326 209 368
rect 263 326 299 368
rect 353 326 389 368
rect 173 310 389 326
rect 173 276 189 310
rect 223 276 257 310
rect 291 276 325 310
rect 359 276 389 310
rect 173 260 389 276
rect 558 330 594 368
rect 648 330 684 368
rect 738 330 774 368
rect 828 330 864 368
rect 920 330 956 368
rect 1010 330 1046 368
rect 558 314 1046 330
rect 558 280 574 314
rect 608 280 642 314
rect 676 280 710 314
rect 744 280 778 314
rect 812 280 846 314
rect 880 280 1046 314
rect 558 264 1046 280
rect 87 222 117 260
rect 173 222 203 260
rect 259 222 289 260
rect 346 222 376 260
rect 558 222 588 264
rect 644 222 674 264
rect 744 222 774 264
rect 830 222 860 264
rect 930 222 960 264
rect 1016 222 1046 264
rect 1102 330 1138 368
rect 1192 330 1228 368
rect 1292 330 1328 368
rect 1382 330 1418 368
rect 1472 330 1508 368
rect 1562 330 1598 368
rect 1652 330 1688 368
rect 1742 330 1778 368
rect 1832 330 1868 368
rect 1922 330 1958 368
rect 2012 330 2048 368
rect 2102 330 2138 368
rect 2192 330 2228 368
rect 2282 330 2318 368
rect 2372 330 2408 368
rect 2472 330 2508 368
rect 1102 314 2508 330
rect 1102 280 1225 314
rect 1259 280 1400 314
rect 1434 280 1580 314
rect 1614 280 1764 314
rect 1798 280 1946 314
rect 1980 280 2135 314
rect 2169 280 2320 314
rect 2354 280 2508 314
rect 1102 264 2508 280
rect 1102 222 1132 264
rect 1188 222 1218 264
rect 1274 222 1304 264
rect 1360 222 1390 264
rect 1446 222 1476 264
rect 1532 222 1562 264
rect 1632 222 1662 264
rect 1718 222 1748 264
rect 1818 222 1848 264
rect 1904 222 1934 264
rect 2004 222 2034 264
rect 2090 222 2120 264
rect 2190 222 2220 264
rect 2276 222 2306 264
rect 2378 222 2408 264
rect 2464 222 2494 264
rect 87 48 117 74
rect 173 48 203 74
rect 259 48 289 74
rect 346 48 376 74
rect 558 48 588 74
rect 644 48 674 74
rect 744 48 774 74
rect 830 48 860 74
rect 930 48 960 74
rect 1016 48 1046 74
rect 1102 48 1132 74
rect 1188 48 1218 74
rect 1274 48 1304 74
rect 1360 48 1390 74
rect 1446 48 1476 74
rect 1532 48 1562 74
rect 1632 48 1662 74
rect 1718 48 1748 74
rect 1818 48 1848 74
rect 1904 48 1934 74
rect 2004 48 2034 74
rect 2090 48 2120 74
rect 2190 48 2220 74
rect 2276 48 2306 74
rect 2378 48 2408 74
rect 2464 48 2494 74
<< polycont >>
rect 51 276 85 310
rect 189 276 223 310
rect 257 276 291 310
rect 325 276 359 310
rect 574 280 608 314
rect 642 280 676 314
rect 710 280 744 314
rect 778 280 812 314
rect 846 280 880 314
rect 1225 280 1259 314
rect 1400 280 1434 314
rect 1580 280 1614 314
rect 1764 280 1798 314
rect 1946 280 1980 314
rect 2135 280 2169 314
rect 2320 280 2354 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 129 580 163 649
rect 129 508 163 546
rect 129 458 163 474
rect 203 580 269 596
rect 203 546 219 580
rect 253 546 269 580
rect 203 497 269 546
rect 203 463 219 497
rect 253 463 269 497
rect 23 406 39 440
rect 73 424 89 440
rect 73 406 169 424
rect 23 390 169 406
rect 25 310 101 356
rect 25 276 51 310
rect 85 276 101 310
rect 25 260 101 276
rect 135 326 169 390
rect 203 414 269 463
rect 309 580 343 649
rect 309 478 343 546
rect 309 428 343 444
rect 383 580 449 596
rect 383 546 399 580
rect 433 546 449 580
rect 383 497 449 546
rect 383 463 399 497
rect 433 463 449 497
rect 203 380 219 414
rect 253 394 269 414
rect 383 414 449 463
rect 383 394 399 414
rect 253 380 399 394
rect 433 380 449 414
rect 203 360 449 380
rect 498 580 548 649
rect 498 546 514 580
rect 498 497 548 546
rect 498 463 514 497
rect 498 414 548 463
rect 498 380 514 414
rect 498 364 548 380
rect 588 580 654 596
rect 588 546 604 580
rect 638 546 654 580
rect 588 497 654 546
rect 588 463 604 497
rect 638 463 654 497
rect 588 414 654 463
rect 694 580 728 649
rect 694 482 728 546
rect 694 432 728 448
rect 768 580 834 596
rect 768 546 784 580
rect 818 546 834 580
rect 768 497 834 546
rect 768 463 784 497
rect 818 463 834 497
rect 588 380 604 414
rect 638 398 654 414
rect 768 414 834 463
rect 874 580 908 649
rect 874 482 908 546
rect 874 432 908 448
rect 950 580 1016 596
rect 950 546 966 580
rect 1000 546 1016 580
rect 950 497 1016 546
rect 950 463 966 497
rect 1000 463 1016 497
rect 768 398 784 414
rect 638 380 784 398
rect 818 398 834 414
rect 950 414 1016 463
rect 950 398 966 414
rect 818 380 966 398
rect 1000 380 1016 414
rect 1056 580 1090 649
rect 1056 503 1090 546
rect 1056 435 1090 469
rect 1056 385 1090 401
rect 1132 580 1198 596
rect 1132 546 1148 580
rect 1182 546 1198 580
rect 1132 497 1198 546
rect 1132 463 1148 497
rect 1182 463 1198 497
rect 1132 424 1198 463
rect 1132 419 1152 424
rect 1132 385 1148 419
rect 1186 390 1198 424
rect 1182 385 1198 390
rect 1232 580 1282 649
rect 1232 546 1248 580
rect 1232 482 1282 546
rect 1232 448 1248 482
rect 1232 385 1282 448
rect 1322 580 1388 596
rect 1322 546 1338 580
rect 1372 546 1388 580
rect 1322 497 1388 546
rect 1322 463 1338 497
rect 1372 463 1388 497
rect 1322 424 1388 463
rect 1322 390 1335 424
rect 1369 418 1388 424
rect 1132 384 1198 385
rect 1322 384 1338 390
rect 1372 384 1388 418
rect 1428 580 1462 649
rect 1428 482 1462 546
rect 1428 385 1462 448
rect 1502 580 1568 596
rect 1502 546 1518 580
rect 1552 546 1568 580
rect 1502 497 1568 546
rect 1502 463 1518 497
rect 1552 463 1568 497
rect 1502 424 1568 463
rect 1502 418 1519 424
rect 1502 384 1518 418
rect 1553 390 1568 424
rect 1552 384 1568 390
rect 1608 580 1642 649
rect 1608 503 1642 546
rect 1608 435 1642 469
rect 1608 385 1642 401
rect 1682 580 1748 596
rect 1682 546 1698 580
rect 1732 546 1748 580
rect 1682 497 1748 546
rect 1682 463 1698 497
rect 1732 463 1748 497
rect 1682 424 1748 463
rect 1682 390 1697 424
rect 1731 418 1748 424
rect 1682 384 1698 390
rect 1732 384 1748 418
rect 1788 580 1822 649
rect 1788 503 1822 546
rect 1788 435 1822 469
rect 1788 385 1822 401
rect 1862 580 1928 596
rect 1862 546 1878 580
rect 1912 546 1928 580
rect 1862 497 1928 546
rect 1862 463 1878 497
rect 1912 463 1928 497
rect 1862 424 1928 463
rect 1862 418 1881 424
rect 1862 384 1878 418
rect 1915 390 1928 424
rect 1912 384 1928 390
rect 1968 580 2002 649
rect 1968 503 2002 546
rect 1968 435 2002 469
rect 1968 385 2002 401
rect 2042 580 2108 596
rect 2042 546 2058 580
rect 2092 546 2108 580
rect 2042 497 2108 546
rect 2042 463 2058 497
rect 2092 463 2108 497
rect 2042 424 2108 463
rect 2042 418 2059 424
rect 2042 384 2058 418
rect 2093 390 2108 424
rect 2092 384 2108 390
rect 2148 580 2182 649
rect 2148 503 2182 546
rect 2148 435 2182 469
rect 2148 385 2182 401
rect 2222 580 2288 596
rect 2222 546 2238 580
rect 2272 546 2288 580
rect 2222 497 2288 546
rect 2222 463 2238 497
rect 2272 463 2288 497
rect 2222 424 2288 463
rect 2222 418 2239 424
rect 2222 384 2238 418
rect 2273 390 2288 424
rect 2272 384 2288 390
rect 2328 580 2378 649
rect 2362 546 2378 580
rect 2328 503 2378 546
rect 2362 469 2378 503
rect 2328 435 2378 469
rect 2362 401 2378 435
rect 2328 385 2378 401
rect 2412 580 2478 596
rect 2412 546 2428 580
rect 2462 546 2478 580
rect 2412 497 2478 546
rect 2412 463 2428 497
rect 2462 463 2478 497
rect 2412 424 2478 463
rect 2412 390 2423 424
rect 2457 414 2478 424
rect 2462 404 2478 414
rect 2518 580 2568 649
rect 2552 546 2568 580
rect 2518 497 2568 546
rect 2552 463 2568 497
rect 2518 414 2568 463
rect 1132 380 1177 384
rect 588 364 1016 380
rect 409 330 449 360
rect 969 351 1016 364
rect 969 350 1081 351
rect 135 310 375 326
rect 135 276 189 310
rect 223 276 257 310
rect 291 276 325 310
rect 359 276 375 310
rect 135 260 375 276
rect 409 314 896 330
rect 409 280 574 314
rect 608 280 642 314
rect 676 280 710 314
rect 744 280 778 314
rect 812 280 846 314
rect 880 280 896 314
rect 409 264 896 280
rect 969 316 1036 350
rect 1070 316 1081 350
rect 969 264 1081 316
rect 135 226 169 260
rect 409 226 443 264
rect 969 230 1021 264
rect 26 210 169 226
rect 26 176 42 210
rect 76 192 169 210
rect 214 210 443 226
rect 26 120 76 176
rect 248 192 387 210
rect 26 86 42 120
rect 26 70 76 86
rect 112 142 178 158
rect 112 108 128 142
rect 162 108 178 142
rect 112 17 178 108
rect 214 120 248 176
rect 371 176 387 192
rect 421 176 443 210
rect 214 70 248 86
rect 284 142 334 158
rect 284 108 300 142
rect 284 17 334 108
rect 371 120 443 176
rect 371 86 387 120
rect 421 86 443 120
rect 371 70 443 86
rect 483 210 549 226
rect 483 176 499 210
rect 533 176 549 210
rect 483 120 549 176
rect 483 86 499 120
rect 533 86 549 120
rect 483 17 549 86
rect 583 210 1021 230
rect 583 176 599 210
rect 633 196 785 210
rect 583 120 633 176
rect 769 176 785 196
rect 819 196 971 210
rect 583 86 599 120
rect 583 70 633 86
rect 669 146 735 162
rect 669 112 685 146
rect 719 112 735 146
rect 669 17 735 112
rect 769 120 819 176
rect 955 176 971 196
rect 1005 196 1021 210
rect 1055 210 1091 226
rect 769 86 785 120
rect 769 70 819 86
rect 855 146 921 162
rect 855 112 871 146
rect 905 112 921 146
rect 855 17 921 112
rect 955 120 1005 176
rect 955 86 971 120
rect 955 70 1005 86
rect 1055 176 1057 210
rect 1055 133 1091 176
rect 1055 99 1057 133
rect 1055 17 1091 99
rect 1127 210 1177 380
rect 1211 316 1225 350
rect 1259 316 1273 350
rect 1322 330 1356 384
rect 1211 314 1273 316
rect 1211 280 1225 314
rect 1259 280 1273 314
rect 1211 264 1273 280
rect 1127 176 1143 210
rect 1127 120 1177 176
rect 1127 86 1143 120
rect 1127 70 1177 86
rect 1213 210 1263 226
rect 1213 176 1229 210
rect 1213 120 1263 176
rect 1213 86 1229 120
rect 1213 17 1263 86
rect 1307 210 1356 330
rect 1390 316 1400 350
rect 1434 316 1443 350
rect 1502 330 1536 384
rect 1390 314 1443 316
rect 1390 280 1400 314
rect 1434 280 1443 314
rect 1390 264 1443 280
rect 1307 176 1315 210
rect 1349 176 1356 210
rect 1307 120 1356 176
rect 1307 86 1315 120
rect 1349 86 1356 120
rect 1307 70 1356 86
rect 1392 210 1435 226
rect 1392 176 1401 210
rect 1392 120 1435 176
rect 1392 86 1401 120
rect 1392 17 1435 86
rect 1477 210 1536 330
rect 1570 316 1580 350
rect 1614 316 1623 350
rect 1682 330 1716 384
rect 1570 314 1623 316
rect 1570 280 1580 314
rect 1614 280 1623 314
rect 1570 264 1623 280
rect 1477 176 1487 210
rect 1521 176 1536 210
rect 1477 120 1536 176
rect 1477 86 1487 120
rect 1521 86 1536 120
rect 1477 70 1536 86
rect 1570 210 1623 226
rect 1570 176 1573 210
rect 1607 176 1623 210
rect 1570 120 1623 176
rect 1570 86 1573 120
rect 1607 86 1623 120
rect 1570 17 1623 86
rect 1657 210 1716 330
rect 1750 316 1764 350
rect 1798 316 1809 350
rect 1862 330 1896 384
rect 1750 314 1809 316
rect 1750 280 1764 314
rect 1798 280 1809 314
rect 1750 264 1809 280
rect 1657 176 1673 210
rect 1707 176 1716 210
rect 1657 120 1716 176
rect 1657 86 1673 120
rect 1707 86 1716 120
rect 1657 70 1716 86
rect 1750 210 1809 226
rect 1750 176 1759 210
rect 1793 176 1809 210
rect 1750 120 1809 176
rect 1750 86 1759 120
rect 1793 86 1809 120
rect 1750 17 1809 86
rect 1843 210 1896 330
rect 1930 316 1946 350
rect 1980 316 1995 350
rect 2042 330 2079 384
rect 1930 314 1995 316
rect 1930 280 1946 314
rect 1980 280 1995 314
rect 1930 264 1995 280
rect 1843 176 1859 210
rect 1893 176 1896 210
rect 1843 120 1896 176
rect 1843 86 1859 120
rect 1893 86 1896 120
rect 1843 70 1896 86
rect 1933 210 1995 226
rect 1933 176 1945 210
rect 1979 176 1995 210
rect 1933 120 1995 176
rect 1933 86 1945 120
rect 1979 86 1995 120
rect 1933 17 1995 86
rect 2029 210 2079 330
rect 2113 316 2135 350
rect 2169 316 2188 350
rect 2113 314 2188 316
rect 2113 280 2135 314
rect 2169 280 2188 314
rect 2113 264 2188 280
rect 2029 176 2045 210
rect 2029 120 2079 176
rect 2029 86 2045 120
rect 2029 70 2079 86
rect 2115 210 2181 226
rect 2115 176 2131 210
rect 2165 176 2181 210
rect 2115 120 2181 176
rect 2115 86 2131 120
rect 2165 86 2181 120
rect 2115 17 2181 86
rect 2222 210 2265 384
rect 2412 380 2428 390
rect 2462 380 2469 404
rect 2299 316 2320 350
rect 2354 316 2378 350
rect 2299 314 2378 316
rect 2299 280 2320 314
rect 2354 280 2378 314
rect 2299 264 2378 280
rect 2412 230 2469 380
rect 2552 380 2568 414
rect 2518 364 2568 380
rect 2222 176 2231 210
rect 2222 120 2265 176
rect 2222 86 2231 120
rect 2222 70 2265 86
rect 2301 210 2367 226
rect 2301 176 2317 210
rect 2351 176 2367 210
rect 2301 120 2367 176
rect 2301 86 2317 120
rect 2351 86 2367 120
rect 2301 17 2367 86
rect 2403 210 2469 230
rect 2403 176 2419 210
rect 2453 176 2469 210
rect 2403 120 2469 176
rect 2403 86 2419 120
rect 2453 86 2469 120
rect 2403 70 2469 86
rect 2503 210 2569 226
rect 2503 176 2519 210
rect 2553 176 2569 210
rect 2503 120 2569 176
rect 2503 86 2519 120
rect 2553 86 2569 120
rect 2503 17 2569 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 1152 419 1186 424
rect 1152 390 1182 419
rect 1182 390 1186 419
rect 1335 418 1369 424
rect 1335 390 1338 418
rect 1338 390 1369 418
rect 1519 418 1553 424
rect 1519 390 1552 418
rect 1552 390 1553 418
rect 1697 418 1731 424
rect 1697 390 1698 418
rect 1698 390 1731 418
rect 1881 418 1915 424
rect 1881 390 1912 418
rect 1912 390 1915 418
rect 2059 418 2093 424
rect 2059 390 2092 418
rect 2092 390 2093 418
rect 2239 418 2273 424
rect 2239 390 2272 418
rect 2272 390 2273 418
rect 2423 414 2457 424
rect 2423 390 2428 414
rect 2428 390 2457 414
rect 1036 316 1070 350
rect 1225 316 1259 350
rect 1400 316 1434 350
rect 1580 316 1614 350
rect 1764 316 1798 350
rect 1946 316 1980 350
rect 2135 316 2169 350
rect 2320 316 2354 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 1140 424 2476 430
rect 1140 390 1152 424
rect 1186 390 1335 424
rect 1369 390 1519 424
rect 1553 390 1697 424
rect 1731 390 1881 424
rect 1915 390 2059 424
rect 2093 390 2239 424
rect 2273 390 2423 424
rect 2457 390 2476 424
rect 1140 384 2476 390
rect 1022 350 2366 356
rect 1022 316 1036 350
rect 1070 316 1225 350
rect 1259 316 1400 350
rect 1434 316 1580 350
rect 1614 316 1764 350
rect 1798 316 1946 350
rect 1980 316 2135 350
rect 2169 316 2320 350
rect 2354 316 2366 350
rect 1022 310 2366 316
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 bufbuf_16
flabel metal1 s 1140 384 2476 430 0 FreeSans 400 0 0 0 X
port 6 nsew
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2592 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3359962
string GDS_START 3339614
<< end >>
