magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 351 2726 704
rect -38 332 527 351
rect 1427 332 2726 351
rect 1629 311 1933 332
<< pwell >>
rect 0 0 2688 49
<< scpmos >>
rect 83 464 119 592
rect 183 464 219 592
rect 267 464 303 592
rect 499 464 535 592
rect 589 464 625 592
rect 703 464 739 592
rect 911 387 947 611
rect 1001 387 1037 611
rect 1209 457 1245 541
rect 1310 461 1346 545
rect 1394 461 1430 545
rect 1519 461 1555 545
rect 1721 347 1757 547
rect 1811 347 1847 547
rect 1960 508 1996 592
rect 2044 508 2080 592
rect 2159 508 2195 592
rect 2249 508 2285 592
rect 2366 424 2402 592
rect 2568 368 2604 592
<< nmoslvt >>
rect 84 88 114 172
rect 282 81 312 165
rect 360 81 390 165
rect 515 81 545 165
rect 593 81 623 165
rect 685 81 715 165
rect 904 119 934 267
rect 1014 119 1044 267
rect 1204 119 1234 203
rect 1290 119 1320 203
rect 1367 119 1397 203
rect 1445 119 1475 203
rect 1629 74 1659 202
rect 1715 74 1745 202
rect 1942 74 1972 158
rect 2014 74 2044 158
rect 2105 74 2135 158
rect 2177 74 2207 158
rect 2376 74 2406 184
rect 2574 74 2604 222
<< ndiff >>
rect 27 147 84 172
rect 27 113 39 147
rect 73 113 84 147
rect 27 88 84 113
rect 114 147 171 172
rect 845 236 904 267
rect 114 113 125 147
rect 159 113 171 147
rect 114 88 171 113
rect 225 127 282 165
rect 225 93 237 127
rect 271 93 282 127
rect 225 81 282 93
rect 312 81 360 165
rect 390 153 515 165
rect 390 119 470 153
rect 504 119 515 153
rect 390 81 515 119
rect 545 81 593 165
rect 623 130 685 165
rect 623 96 636 130
rect 670 96 685 130
rect 623 81 685 96
rect 715 130 772 165
rect 715 96 726 130
rect 760 96 772 130
rect 715 81 772 96
rect 835 150 904 236
rect 835 116 847 150
rect 881 119 904 150
rect 934 150 1014 267
rect 934 119 957 150
rect 881 116 889 119
rect 835 93 889 116
rect 949 116 957 119
rect 991 119 1014 150
rect 1044 235 1097 267
rect 1044 201 1055 235
rect 1089 201 1097 235
rect 1044 165 1097 201
rect 1044 131 1055 165
rect 1089 131 1097 165
rect 1044 119 1097 131
rect 1151 179 1204 203
rect 1151 145 1159 179
rect 1193 145 1204 179
rect 1151 119 1204 145
rect 1234 179 1290 203
rect 1234 145 1245 179
rect 1279 145 1290 179
rect 1234 119 1290 145
rect 1320 119 1367 203
rect 1397 119 1445 203
rect 1475 202 1599 203
rect 1475 119 1629 202
rect 991 116 999 119
rect 949 93 999 116
rect 1490 82 1629 119
rect 1490 48 1502 82
rect 1536 74 1629 82
rect 1659 179 1715 202
rect 1659 145 1670 179
rect 1704 145 1715 179
rect 1659 74 1715 145
rect 1745 158 1795 202
rect 2517 210 2574 222
rect 1745 129 1942 158
rect 1745 95 1897 129
rect 1931 95 1942 129
rect 1745 74 1942 95
rect 1972 74 2014 158
rect 2044 133 2105 158
rect 2044 99 2055 133
rect 2089 99 2105 133
rect 2044 74 2105 99
rect 2135 74 2177 158
rect 2207 133 2264 158
rect 2207 99 2218 133
rect 2252 99 2264 133
rect 2207 74 2264 99
rect 2318 117 2376 184
rect 2318 83 2330 117
rect 2364 83 2376 117
rect 2318 74 2376 83
rect 2406 146 2463 184
rect 2406 112 2417 146
rect 2451 112 2463 146
rect 2406 74 2463 112
rect 2517 176 2529 210
rect 2563 176 2574 210
rect 2517 120 2574 176
rect 2517 86 2529 120
rect 2563 86 2574 120
rect 2517 74 2574 86
rect 2604 210 2661 222
rect 2604 176 2615 210
rect 2649 176 2661 210
rect 2604 120 2661 176
rect 2604 86 2615 120
rect 2649 86 2661 120
rect 2604 74 2661 86
rect 1536 48 1548 74
rect 1490 36 1548 48
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 464 83 476
rect 119 580 183 592
rect 119 546 139 580
rect 173 546 183 580
rect 119 510 183 546
rect 119 476 139 510
rect 173 476 183 510
rect 119 464 183 476
rect 219 464 267 592
rect 303 580 499 592
rect 303 546 313 580
rect 347 546 384 580
rect 418 546 454 580
rect 488 546 499 580
rect 303 510 499 546
rect 303 476 313 510
rect 347 476 384 510
rect 418 476 454 510
rect 488 476 499 510
rect 303 464 499 476
rect 535 464 589 592
rect 625 575 703 592
rect 625 541 635 575
rect 669 541 703 575
rect 625 464 703 541
rect 739 580 795 592
rect 739 546 749 580
rect 783 546 795 580
rect 739 512 795 546
rect 739 478 749 512
rect 783 478 795 512
rect 739 464 795 478
rect 855 441 911 611
rect 855 407 867 441
rect 901 407 911 441
rect 855 387 911 407
rect 947 594 1001 611
rect 947 560 957 594
rect 991 560 1001 594
rect 947 387 1001 560
rect 1037 441 1093 611
rect 1037 407 1047 441
rect 1081 407 1093 441
rect 1037 387 1093 407
rect 1445 582 1504 594
rect 1445 548 1457 582
rect 1491 548 1504 582
rect 1445 545 1504 548
rect 1862 560 1960 592
rect 1862 547 1895 560
rect 1260 541 1310 545
rect 1153 516 1209 541
rect 1153 482 1165 516
rect 1199 482 1209 516
rect 1153 457 1209 482
rect 1245 528 1310 541
rect 1245 494 1266 528
rect 1300 494 1310 528
rect 1245 461 1310 494
rect 1346 461 1394 545
rect 1430 461 1519 545
rect 1555 523 1611 545
rect 1555 489 1565 523
rect 1599 489 1611 523
rect 1555 461 1611 489
rect 1665 535 1721 547
rect 1665 501 1677 535
rect 1711 501 1721 535
rect 1665 467 1721 501
rect 1245 457 1295 461
rect 1665 433 1677 467
rect 1711 433 1721 467
rect 1665 399 1721 433
rect 1665 365 1677 399
rect 1711 365 1721 399
rect 1665 347 1721 365
rect 1757 535 1811 547
rect 1757 501 1767 535
rect 1801 501 1811 535
rect 1757 464 1811 501
rect 1757 430 1767 464
rect 1801 430 1811 464
rect 1757 393 1811 430
rect 1757 359 1767 393
rect 1801 359 1811 393
rect 1757 347 1811 359
rect 1847 526 1895 547
rect 1929 526 1960 560
rect 1847 508 1960 526
rect 1996 508 2044 592
rect 2080 567 2159 592
rect 2080 533 2097 567
rect 2131 533 2159 567
rect 2080 508 2159 533
rect 2195 567 2249 592
rect 2195 533 2205 567
rect 2239 533 2249 567
rect 2195 508 2249 533
rect 2285 580 2366 592
rect 2285 546 2312 580
rect 2346 546 2366 580
rect 2285 508 2366 546
rect 1847 347 1897 508
rect 2300 470 2366 508
rect 2300 436 2312 470
rect 2346 436 2366 470
rect 2300 424 2366 436
rect 2402 580 2458 592
rect 2402 546 2412 580
rect 2446 546 2458 580
rect 2402 470 2458 546
rect 2402 436 2412 470
rect 2446 436 2458 470
rect 2402 424 2458 436
rect 2512 580 2568 592
rect 2512 546 2524 580
rect 2558 546 2568 580
rect 2512 497 2568 546
rect 2512 463 2524 497
rect 2558 463 2568 497
rect 2512 414 2568 463
rect 2512 380 2524 414
rect 2558 380 2568 414
rect 2512 368 2568 380
rect 2604 580 2660 592
rect 2604 546 2614 580
rect 2648 546 2660 580
rect 2604 497 2660 546
rect 2604 463 2614 497
rect 2648 463 2660 497
rect 2604 414 2660 463
rect 2604 380 2614 414
rect 2648 380 2660 414
rect 2604 368 2660 380
<< ndiffc >>
rect 39 113 73 147
rect 125 113 159 147
rect 237 93 271 127
rect 470 119 504 153
rect 636 96 670 130
rect 726 96 760 130
rect 847 116 881 150
rect 957 116 991 150
rect 1055 201 1089 235
rect 1055 131 1089 165
rect 1159 145 1193 179
rect 1245 145 1279 179
rect 1502 48 1536 82
rect 1670 145 1704 179
rect 1897 95 1931 129
rect 2055 99 2089 133
rect 2218 99 2252 133
rect 2330 83 2364 117
rect 2417 112 2451 146
rect 2529 176 2563 210
rect 2529 86 2563 120
rect 2615 176 2649 210
rect 2615 86 2649 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 139 546 173 580
rect 139 476 173 510
rect 313 546 347 580
rect 384 546 418 580
rect 454 546 488 580
rect 313 476 347 510
rect 384 476 418 510
rect 454 476 488 510
rect 635 541 669 575
rect 749 546 783 580
rect 749 478 783 512
rect 867 407 901 441
rect 957 560 991 594
rect 1047 407 1081 441
rect 1457 548 1491 582
rect 1165 482 1199 516
rect 1266 494 1300 528
rect 1565 489 1599 523
rect 1677 501 1711 535
rect 1677 433 1711 467
rect 1677 365 1711 399
rect 1767 501 1801 535
rect 1767 430 1801 464
rect 1767 359 1801 393
rect 1895 526 1929 560
rect 2097 533 2131 567
rect 2205 533 2239 567
rect 2312 546 2346 580
rect 2312 436 2346 470
rect 2412 546 2446 580
rect 2412 436 2446 470
rect 2524 546 2558 580
rect 2524 463 2558 497
rect 2524 380 2558 414
rect 2614 546 2648 580
rect 2614 463 2648 497
rect 2614 380 2648 414
<< poly >>
rect 83 592 119 618
rect 183 592 219 618
rect 267 592 303 618
rect 499 592 535 618
rect 589 592 625 618
rect 703 592 739 618
rect 911 611 947 643
rect 1001 611 1037 643
rect 1108 615 1847 645
rect 83 367 119 464
rect 183 367 219 464
rect 267 445 303 464
rect 267 415 353 445
rect 499 432 535 464
rect 589 449 625 464
rect 703 449 739 464
rect 83 351 225 367
rect 83 337 107 351
rect 84 317 107 337
rect 141 317 175 351
rect 209 317 225 351
rect 84 301 225 317
rect 323 318 353 415
rect 401 416 535 432
rect 401 382 417 416
rect 451 382 485 416
rect 519 382 535 416
rect 401 366 535 382
rect 577 406 643 449
rect 577 372 593 406
rect 627 372 643 406
rect 577 338 643 372
rect 84 172 114 301
rect 323 288 384 318
rect 354 253 384 288
rect 469 302 535 318
rect 469 268 485 302
rect 519 268 535 302
rect 577 304 593 338
rect 627 304 643 338
rect 577 288 643 304
rect 685 432 739 449
rect 685 416 823 432
rect 685 382 773 416
rect 807 382 823 416
rect 685 370 823 382
rect 911 372 947 387
rect 685 366 819 370
rect 209 237 275 253
rect 209 203 225 237
rect 259 217 275 237
rect 354 237 420 253
rect 469 252 535 268
rect 259 203 312 217
rect 209 187 312 203
rect 354 203 370 237
rect 404 203 420 237
rect 354 187 420 203
rect 505 210 535 252
rect 282 165 312 187
rect 360 165 390 187
rect 505 180 545 210
rect 515 165 545 180
rect 593 165 623 288
rect 685 165 715 366
rect 866 351 947 372
rect 1001 370 1037 387
rect 1108 370 1138 615
rect 1209 541 1245 567
rect 1310 545 1346 615
rect 1394 545 1430 571
rect 1519 545 1555 571
rect 1721 547 1757 573
rect 1811 547 1847 615
rect 1960 592 1996 618
rect 2044 592 2080 618
rect 2159 592 2195 618
rect 2249 592 2285 618
rect 2366 592 2402 618
rect 2568 592 2604 618
rect 1209 375 1245 457
rect 1310 435 1346 461
rect 862 339 947 351
rect 862 324 878 339
rect 757 308 878 324
rect 757 274 773 308
rect 807 305 878 308
rect 912 318 947 339
rect 990 339 1138 370
rect 912 305 944 318
rect 807 282 944 305
rect 990 305 1006 339
rect 1040 305 1138 339
rect 1180 359 1246 375
rect 1394 361 1430 461
rect 1519 429 1555 461
rect 1519 413 1633 429
rect 1519 379 1583 413
rect 1617 379 1633 413
rect 1519 363 1633 379
rect 1180 325 1196 359
rect 1230 345 1246 359
rect 1367 345 1470 361
rect 1230 325 1320 345
rect 1180 315 1320 325
rect 1180 309 1246 315
rect 990 297 1138 305
rect 990 296 1139 297
rect 990 293 1140 296
rect 990 290 1141 293
rect 990 282 1142 290
rect 807 274 823 282
rect 757 258 823 274
rect 904 267 934 282
rect 1014 267 1044 282
rect 1112 267 1142 282
rect 84 62 114 88
rect 904 93 934 119
rect 1112 237 1234 267
rect 1204 203 1234 237
rect 1290 203 1320 315
rect 1367 311 1420 345
rect 1454 311 1470 345
rect 1367 295 1470 311
rect 1367 203 1397 295
rect 1519 253 1549 363
rect 1960 476 1996 508
rect 1929 460 1996 476
rect 1929 426 1945 460
rect 1979 426 1996 460
rect 1929 410 1996 426
rect 2044 368 2080 508
rect 2159 430 2195 508
rect 1721 319 1757 347
rect 1633 315 1757 319
rect 1445 223 1549 253
rect 1597 299 1757 315
rect 1811 332 1847 347
rect 2033 338 2080 368
rect 2128 414 2195 430
rect 2128 380 2144 414
rect 2178 380 2195 414
rect 2128 364 2195 380
rect 2249 398 2285 508
rect 2366 398 2402 424
rect 2249 368 2402 398
rect 1811 302 1955 332
rect 1597 265 1613 299
rect 1647 289 1757 299
rect 1647 265 1663 289
rect 1597 249 1663 265
rect 1445 203 1475 223
rect 1629 202 1659 249
rect 1817 247 1883 254
rect 1715 238 1883 247
rect 1715 217 1833 238
rect 1715 202 1745 217
rect 1817 204 1833 217
rect 1867 204 1883 238
rect 1014 93 1044 119
rect 1204 93 1234 119
rect 1290 93 1320 119
rect 1367 93 1397 119
rect 282 55 312 81
rect 360 55 390 81
rect 515 55 545 81
rect 593 55 623 81
rect 685 51 715 81
rect 1445 51 1475 119
rect 685 21 1475 51
rect 1817 188 1883 204
rect 1925 224 1955 302
rect 1997 322 2063 338
rect 1997 288 2013 322
rect 2047 288 2063 322
rect 2128 290 2158 364
rect 1997 272 2063 288
rect 1925 194 1972 224
rect 1942 158 1972 194
rect 2014 158 2044 272
rect 2105 260 2158 290
rect 2249 270 2279 368
rect 2568 326 2604 368
rect 2448 310 2604 326
rect 2448 276 2464 310
rect 2498 276 2532 310
rect 2566 276 2604 310
rect 2105 158 2135 260
rect 2213 254 2406 270
rect 2448 260 2604 276
rect 2213 220 2229 254
rect 2263 240 2406 254
rect 2263 220 2279 240
rect 2213 218 2279 220
rect 2177 188 2279 218
rect 2177 158 2207 188
rect 2376 184 2406 240
rect 2574 222 2604 260
rect 1629 48 1659 74
rect 1715 48 1745 74
rect 1942 48 1972 74
rect 2014 48 2044 74
rect 2105 48 2135 74
rect 2177 48 2207 74
rect 2376 48 2406 74
rect 2574 48 2604 74
<< polycont >>
rect 107 317 141 351
rect 175 317 209 351
rect 417 382 451 416
rect 485 382 519 416
rect 593 372 627 406
rect 485 268 519 302
rect 593 304 627 338
rect 773 382 807 416
rect 225 203 259 237
rect 370 203 404 237
rect 773 274 807 308
rect 878 305 912 339
rect 1006 305 1040 339
rect 1583 379 1617 413
rect 1196 325 1230 359
rect 1420 311 1454 345
rect 1945 426 1979 460
rect 2144 380 2178 414
rect 1613 265 1647 299
rect 1833 204 1867 238
rect 2013 288 2047 322
rect 2464 276 2498 310
rect 2532 276 2566 310
rect 2229 220 2263 254
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 435 89 476
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 510 189 546
rect 123 476 139 510
rect 173 476 189 510
rect 123 469 189 476
rect 297 580 511 596
rect 297 546 313 580
rect 347 546 384 580
rect 418 546 454 580
rect 488 546 511 580
rect 297 510 511 546
rect 619 575 685 649
rect 619 541 635 575
rect 669 541 685 575
rect 619 537 685 541
rect 733 580 799 596
rect 733 546 749 580
rect 783 546 799 580
rect 941 594 1007 649
rect 941 560 957 594
rect 991 560 1007 594
rect 1441 582 1508 649
rect 297 476 313 510
rect 347 476 384 510
rect 418 476 454 510
rect 488 503 511 510
rect 733 526 799 546
rect 1441 548 1457 582
rect 1491 548 1508 582
rect 1165 526 1215 545
rect 733 516 1215 526
rect 733 512 1165 516
rect 733 503 749 512
rect 488 478 749 503
rect 783 491 1165 512
rect 783 478 799 491
rect 1199 482 1215 516
rect 488 476 757 478
rect 297 469 757 476
rect 689 466 757 469
rect 23 416 541 435
rect 23 401 417 416
rect 23 253 57 401
rect 407 382 417 401
rect 451 382 485 416
rect 519 382 541 416
rect 91 351 359 367
rect 407 366 541 382
rect 589 406 655 430
rect 589 372 593 406
rect 627 372 655 406
rect 91 317 107 351
rect 141 317 175 351
rect 209 332 359 351
rect 589 338 655 372
rect 209 317 545 332
rect 91 302 545 317
rect 91 298 485 302
rect 469 268 485 298
rect 519 268 545 302
rect 589 304 593 338
rect 627 304 655 338
rect 589 288 655 304
rect 23 237 275 253
rect 23 210 225 237
rect 23 147 73 210
rect 209 203 225 210
rect 259 203 275 237
rect 209 187 275 203
rect 313 237 420 253
rect 469 252 545 268
rect 313 203 370 237
rect 404 203 420 237
rect 689 218 723 466
rect 784 432 833 444
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 867 441 917 457
rect 901 434 917 441
rect 1031 441 1126 457
rect 901 407 996 434
rect 867 390 996 407
rect 1031 407 1047 441
rect 1081 407 1126 441
rect 1165 443 1215 482
rect 1250 528 1376 545
rect 1441 532 1508 548
rect 1250 494 1266 528
rect 1300 498 1376 528
rect 1549 523 1615 549
rect 1549 498 1565 523
rect 1300 494 1565 498
rect 1250 489 1565 494
rect 1599 489 1615 523
rect 1250 477 1615 489
rect 1342 464 1615 477
rect 1677 535 1711 649
rect 1858 560 2063 576
rect 1677 467 1711 501
rect 1165 409 1308 443
rect 1031 394 1126 407
rect 807 382 833 390
rect 757 366 833 382
rect 962 360 996 390
rect 1090 375 1126 394
rect 867 339 928 355
rect 867 332 878 339
rect 23 113 39 147
rect 23 84 73 113
rect 109 147 175 176
rect 313 162 420 203
rect 454 184 723 218
rect 757 308 878 332
rect 757 274 773 308
rect 807 305 878 308
rect 912 305 928 339
rect 807 274 928 305
rect 757 252 928 274
rect 962 339 1056 360
rect 962 305 1006 339
rect 1040 305 1056 339
rect 962 289 1056 305
rect 1090 359 1240 375
rect 1090 325 1196 359
rect 1230 325 1240 359
rect 1090 309 1240 325
rect 757 184 839 252
rect 962 218 1009 289
rect 1090 253 1126 309
rect 1274 274 1308 409
rect 873 184 1009 218
rect 1043 235 1126 253
rect 1043 201 1055 235
rect 1089 222 1126 235
rect 1160 240 1308 274
rect 1089 201 1124 222
rect 1160 207 1195 240
rect 109 113 125 147
rect 159 113 175 147
rect 454 153 520 184
rect 109 17 175 113
rect 221 127 287 128
rect 221 93 237 127
rect 271 93 287 127
rect 454 119 470 153
rect 504 119 520 153
rect 873 150 907 184
rect 1043 165 1124 201
rect 612 130 682 150
rect 221 85 287 93
rect 612 96 636 130
rect 670 96 682 130
rect 612 85 682 96
rect 221 51 682 85
rect 718 130 776 150
rect 718 96 726 130
rect 760 96 776 130
rect 827 116 847 150
rect 881 116 907 150
rect 827 100 907 116
rect 941 116 957 150
rect 991 116 1007 150
rect 718 17 776 96
rect 941 17 1007 116
rect 1043 131 1055 165
rect 1089 131 1124 165
rect 1043 85 1124 131
rect 1159 179 1195 207
rect 1342 206 1376 464
rect 1193 145 1195 179
rect 1159 119 1195 145
rect 1229 179 1376 206
rect 1410 345 1465 361
rect 1410 311 1420 345
rect 1454 311 1465 345
rect 1410 218 1465 311
rect 1499 315 1533 464
rect 1567 424 1633 430
rect 1601 413 1633 424
rect 1567 379 1583 390
rect 1617 379 1633 413
rect 1567 363 1633 379
rect 1677 399 1711 433
rect 1677 349 1711 365
rect 1745 535 1801 551
rect 1745 501 1767 535
rect 1858 526 1895 560
rect 1929 526 2063 560
rect 1858 510 2063 526
rect 1745 464 1801 501
rect 1745 430 1767 464
rect 1745 393 1801 430
rect 1745 359 1767 393
rect 1745 343 1801 359
rect 1849 460 1995 476
rect 1849 426 1945 460
rect 1979 426 1995 460
rect 1849 425 1995 426
rect 1499 299 1663 315
rect 1499 265 1613 299
rect 1647 265 1663 299
rect 1499 252 1663 265
rect 1745 218 1779 343
rect 1849 254 1883 425
rect 2029 391 2063 510
rect 2097 567 2147 649
rect 2131 533 2147 567
rect 2097 504 2147 533
rect 2189 567 2262 596
rect 2189 533 2205 567
rect 2239 533 2262 567
rect 2189 504 2262 533
rect 1410 184 1779 218
rect 1813 238 1883 254
rect 1813 204 1833 238
rect 1867 204 1883 238
rect 1813 188 1883 204
rect 1917 357 2063 391
rect 2128 424 2194 430
rect 2128 390 2143 424
rect 2177 414 2194 424
rect 2128 380 2144 390
rect 2178 380 2194 414
rect 2128 364 2194 380
rect 1917 253 1951 357
rect 2228 323 2262 504
rect 2296 580 2362 649
rect 2296 546 2312 580
rect 2346 546 2362 580
rect 2296 470 2362 546
rect 2296 436 2312 470
rect 2346 436 2362 470
rect 2296 420 2362 436
rect 2396 580 2462 596
rect 2396 546 2412 580
rect 2446 546 2462 580
rect 2396 470 2462 546
rect 2396 436 2412 470
rect 2446 436 2462 470
rect 2396 420 2462 436
rect 2417 326 2462 420
rect 2508 580 2574 649
rect 2508 546 2524 580
rect 2558 546 2574 580
rect 2508 497 2574 546
rect 2508 463 2524 497
rect 2558 463 2574 497
rect 2508 414 2574 463
rect 2508 380 2524 414
rect 2558 380 2574 414
rect 2508 364 2574 380
rect 2614 580 2665 596
rect 2648 546 2665 580
rect 2614 497 2665 546
rect 2648 463 2665 497
rect 2614 414 2665 463
rect 2648 380 2665 414
rect 1997 322 2347 323
rect 1997 288 2013 322
rect 2047 289 2347 322
rect 2047 288 2063 289
rect 1997 287 2063 288
rect 2213 254 2279 255
rect 2213 253 2229 254
rect 1917 220 2229 253
rect 2263 220 2279 254
rect 1917 219 2279 220
rect 1229 145 1245 179
rect 1279 172 1376 179
rect 1654 179 1731 184
rect 1279 145 1294 172
rect 1229 119 1294 145
rect 1410 116 1620 150
rect 1654 145 1670 179
rect 1704 145 1731 179
rect 1654 119 1731 145
rect 1410 85 1444 116
rect 1043 51 1444 85
rect 1586 85 1620 116
rect 1813 85 1847 188
rect 1917 154 1951 219
rect 2313 185 2347 289
rect 1486 48 1502 82
rect 1536 48 1552 82
rect 1586 51 1847 85
rect 1881 129 1951 154
rect 1881 95 1897 129
rect 1931 95 1951 129
rect 1881 70 1951 95
rect 2039 133 2105 162
rect 2039 99 2055 133
rect 2089 99 2105 133
rect 1486 17 1552 48
rect 2039 17 2105 99
rect 2202 151 2347 185
rect 2417 310 2574 326
rect 2417 276 2464 310
rect 2498 276 2532 310
rect 2566 276 2574 310
rect 2417 260 2574 276
rect 2202 133 2268 151
rect 2202 99 2218 133
rect 2252 99 2268 133
rect 2417 146 2467 260
rect 2614 226 2665 380
rect 2202 70 2268 99
rect 2314 83 2330 117
rect 2364 83 2381 117
rect 2314 17 2381 83
rect 2451 112 2467 146
rect 2417 70 2467 112
rect 2513 210 2563 226
rect 2513 176 2529 210
rect 2513 120 2563 176
rect 2513 86 2529 120
rect 2513 17 2563 86
rect 2599 210 2665 226
rect 2599 176 2615 210
rect 2649 176 2665 210
rect 2599 120 2665 176
rect 2599 86 2615 120
rect 2649 86 2665 120
rect 2599 70 2665 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1567 413 1601 424
rect 1567 390 1583 413
rect 1583 390 1601 413
rect 2143 414 2177 424
rect 2143 390 2144 414
rect 2144 390 2177 414
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfrtp_1
flabel comment s 1507 630 1507 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1094 36 1094 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 2143 390 2177 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2623 94 2657 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2688 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 231846
string GDS_START 210444
<< end >>
