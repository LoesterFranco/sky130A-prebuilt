magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 98 153 166 335
rect 200 153 276 285
rect 399 289 1267 345
rect 1221 171 1267 289
rect 899 123 1267 171
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 353 69 493
rect 103 369 196 527
rect 240 353 291 493
rect 333 421 382 493
rect 416 455 492 527
rect 536 421 570 493
rect 614 455 680 527
rect 724 421 1257 493
rect 333 387 1257 421
rect 399 379 1257 387
rect 17 255 64 353
rect 17 221 30 255
rect 17 133 64 221
rect 240 319 365 353
rect 310 255 365 319
rect 310 205 832 255
rect 866 221 942 255
rect 976 221 1187 255
rect 866 205 1187 221
rect 17 56 69 133
rect 310 119 365 205
rect 103 17 196 119
rect 240 51 365 119
rect 399 131 865 171
rect 399 51 465 131
rect 499 17 575 97
rect 619 55 653 131
rect 687 17 763 97
rect 807 89 865 131
rect 807 51 1257 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 30 221 64 255
rect 942 221 976 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< obsm1 >>
rect 17 255 988 261
rect 17 221 30 255
rect 64 233 942 255
rect 64 221 76 233
rect 17 215 76 221
rect 930 221 942 233
rect 976 221 988 255
rect 930 215 988 221
<< labels >>
rlabel locali s 98 153 166 335 6 A
port 1 nsew signal input
rlabel locali s 200 153 276 285 6 TE_B
port 2 nsew signal input
rlabel locali s 1221 171 1267 289 6 Z
port 3 nsew signal output
rlabel locali s 899 123 1267 171 6 Z
port 3 nsew signal output
rlabel locali s 399 289 1267 345 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1990636
string GDS_START 1980902
<< end >>
