magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 281 47 311 177
rect 375 47 405 177
rect 469 47 499 177
rect 674 47 704 177
rect 768 47 798 177
rect 862 47 892 177
rect 956 47 986 177
<< pmoshvt >>
rect 81 297 117 497
rect 289 309 325 497
rect 383 309 419 497
rect 477 309 513 497
rect 571 309 607 497
rect 676 297 712 497
rect 770 297 806 497
rect 864 297 900 497
rect 958 297 994 497
<< ndiff >>
rect 27 106 89 177
rect 27 72 35 106
rect 69 72 89 106
rect 27 47 89 72
rect 119 89 183 177
rect 119 55 129 89
rect 163 55 183 89
rect 119 47 183 55
rect 213 124 281 177
rect 213 90 227 124
rect 261 90 281 124
rect 213 47 281 90
rect 311 89 375 177
rect 311 55 321 89
rect 355 55 375 89
rect 311 47 375 55
rect 405 124 469 177
rect 405 90 415 124
rect 449 90 469 124
rect 405 47 469 90
rect 499 89 555 177
rect 499 55 509 89
rect 543 55 555 89
rect 499 47 555 55
rect 622 124 674 177
rect 622 90 630 124
rect 664 90 674 124
rect 622 47 674 90
rect 704 169 768 177
rect 704 135 724 169
rect 758 135 768 169
rect 704 47 768 135
rect 798 89 862 177
rect 798 55 818 89
rect 852 55 862 89
rect 798 47 862 55
rect 892 169 956 177
rect 892 135 912 169
rect 946 135 956 169
rect 892 47 956 135
rect 986 89 1052 177
rect 986 55 1006 89
rect 1040 55 1052 89
rect 986 47 1052 55
<< pdiff >>
rect 27 450 81 497
rect 27 416 35 450
rect 69 416 81 450
rect 27 297 81 416
rect 117 485 171 497
rect 117 451 129 485
rect 163 451 171 485
rect 117 297 171 451
rect 235 465 289 497
rect 235 431 243 465
rect 277 431 289 465
rect 235 309 289 431
rect 325 489 383 497
rect 325 455 337 489
rect 371 455 383 489
rect 325 421 383 455
rect 325 387 337 421
rect 371 387 383 421
rect 325 309 383 387
rect 419 477 477 497
rect 419 443 431 477
rect 465 443 477 477
rect 419 409 477 443
rect 419 375 431 409
rect 465 375 477 409
rect 419 309 477 375
rect 513 489 571 497
rect 513 455 525 489
rect 559 455 571 489
rect 513 421 571 455
rect 513 387 525 421
rect 559 387 571 421
rect 513 309 571 387
rect 607 477 676 497
rect 607 443 625 477
rect 659 443 676 477
rect 607 409 676 443
rect 607 375 625 409
rect 659 375 676 409
rect 607 309 676 375
rect 624 297 676 309
rect 712 407 770 497
rect 712 373 724 407
rect 758 373 770 407
rect 712 339 770 373
rect 712 305 724 339
rect 758 305 770 339
rect 712 297 770 305
rect 806 477 864 497
rect 806 443 818 477
rect 852 443 864 477
rect 806 409 864 443
rect 806 375 818 409
rect 852 375 864 409
rect 806 297 864 375
rect 900 407 958 497
rect 900 373 912 407
rect 946 373 958 407
rect 900 339 958 373
rect 900 305 912 339
rect 946 305 958 339
rect 900 297 958 305
rect 994 477 1048 497
rect 994 443 1006 477
rect 1040 443 1048 477
rect 994 409 1048 443
rect 994 375 1006 409
rect 1040 375 1048 409
rect 994 297 1048 375
<< ndiffc >>
rect 35 72 69 106
rect 129 55 163 89
rect 227 90 261 124
rect 321 55 355 89
rect 415 90 449 124
rect 509 55 543 89
rect 630 90 664 124
rect 724 135 758 169
rect 818 55 852 89
rect 912 135 946 169
rect 1006 55 1040 89
<< pdiffc >>
rect 35 416 69 450
rect 129 451 163 485
rect 243 431 277 465
rect 337 455 371 489
rect 337 387 371 421
rect 431 443 465 477
rect 431 375 465 409
rect 525 455 559 489
rect 525 387 559 421
rect 625 443 659 477
rect 625 375 659 409
rect 724 373 758 407
rect 724 305 758 339
rect 818 443 852 477
rect 818 375 852 409
rect 912 373 946 407
rect 912 305 946 339
rect 1006 443 1040 477
rect 1006 375 1040 409
<< poly >>
rect 81 497 117 523
rect 289 497 325 523
rect 383 497 419 523
rect 477 497 513 523
rect 571 497 607 523
rect 676 497 712 523
rect 770 497 806 523
rect 864 497 900 523
rect 958 497 994 523
rect 81 282 117 297
rect 289 294 325 309
rect 383 294 419 309
rect 477 294 513 309
rect 571 294 607 309
rect 79 265 119 282
rect 21 249 119 265
rect 287 264 609 294
rect 676 282 712 297
rect 770 282 806 297
rect 864 282 900 297
rect 958 282 994 297
rect 21 215 32 249
rect 66 222 119 249
rect 545 249 609 264
rect 66 215 499 222
rect 21 199 499 215
rect 545 215 555 249
rect 589 215 609 249
rect 545 199 609 215
rect 674 265 714 282
rect 768 265 808 282
rect 674 259 808 265
rect 862 259 902 282
rect 956 261 996 282
rect 956 259 1050 261
rect 674 249 1050 259
rect 674 215 858 249
rect 892 215 932 249
rect 966 215 1000 249
rect 1034 215 1050 249
rect 674 205 1050 215
rect 674 199 798 205
rect 89 192 499 199
rect 89 177 119 192
rect 183 177 213 192
rect 281 177 311 192
rect 375 177 405 192
rect 469 177 499 192
rect 674 177 704 199
rect 768 177 798 199
rect 862 177 892 205
rect 956 203 1050 205
rect 956 177 986 203
rect 89 21 119 47
rect 183 21 213 47
rect 281 21 311 47
rect 375 21 405 47
rect 469 21 499 47
rect 674 21 704 47
rect 768 21 798 47
rect 862 21 892 47
rect 956 21 986 47
<< polycont >>
rect 32 215 66 249
rect 555 215 589 249
rect 858 215 892 249
rect 932 215 966 249
rect 1000 215 1034 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 450 69 493
rect 17 416 35 450
rect 103 485 185 527
rect 103 451 129 485
rect 163 451 185 485
rect 103 425 185 451
rect 235 465 277 493
rect 235 431 243 465
rect 17 391 69 416
rect 17 357 185 391
rect 17 249 66 323
rect 17 215 32 249
rect 17 199 66 215
rect 100 265 185 357
rect 235 345 277 431
rect 321 489 387 527
rect 321 455 337 489
rect 371 455 387 489
rect 321 421 387 455
rect 321 387 337 421
rect 371 387 387 421
rect 321 379 387 387
rect 431 477 465 493
rect 431 409 465 443
rect 509 489 581 527
rect 509 455 525 489
rect 559 455 581 489
rect 509 421 581 455
rect 509 387 525 421
rect 559 387 581 421
rect 509 379 581 387
rect 625 477 1082 493
rect 659 459 818 477
rect 625 409 659 443
rect 852 459 1006 477
rect 431 345 465 375
rect 625 345 659 375
rect 235 311 659 345
rect 698 407 774 425
rect 698 373 724 407
rect 758 373 774 407
rect 698 339 774 373
rect 818 409 852 443
rect 1040 443 1082 477
rect 818 357 852 375
rect 886 407 962 425
rect 886 373 912 407
rect 946 373 962 407
rect 698 305 724 339
rect 758 323 774 339
rect 886 339 962 373
rect 886 323 912 339
rect 758 305 912 323
rect 946 305 962 339
rect 698 289 962 305
rect 1006 409 1082 443
rect 1040 375 1082 409
rect 1006 289 1082 375
rect 100 249 664 265
rect 100 215 555 249
rect 589 215 664 249
rect 100 199 664 215
rect 100 165 149 199
rect 698 170 806 289
rect 842 249 1082 255
rect 842 215 858 249
rect 892 215 932 249
rect 966 215 1000 249
rect 1034 215 1082 249
rect 842 204 1082 215
rect 698 169 1082 170
rect 17 131 149 165
rect 227 131 664 165
rect 17 106 69 131
rect 17 72 35 106
rect 227 124 261 131
rect 17 51 69 72
rect 103 89 179 97
rect 103 55 129 89
rect 163 55 179 89
rect 103 17 179 55
rect 415 124 449 131
rect 227 51 261 90
rect 295 89 371 97
rect 295 55 321 89
rect 355 55 371 89
rect 295 17 371 55
rect 597 124 664 131
rect 698 135 724 169
rect 758 135 912 169
rect 946 135 1082 169
rect 698 127 1082 135
rect 415 51 449 90
rect 483 89 561 97
rect 483 55 509 89
rect 543 55 561 89
rect 483 17 561 55
rect 597 90 630 124
rect 664 90 1082 93
rect 597 89 1082 90
rect 597 55 818 89
rect 852 55 1006 89
rect 1040 55 1082 89
rect 597 51 1082 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 TE
port 2 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 TE
port 2 nsew
flabel corelocali s 950 221 984 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 850 221 884 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1039 221 1073 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 850 289 884 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 748 289 782 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 748 153 782 187 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 748 221 782 255 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
rlabel comment s 0 0 0 0 4 einvp_4
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2057858
string GDS_START 2049542
<< end >>
