magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2392 561
rect 103 427 169 527
rect 17 195 87 325
rect 286 427 357 527
rect 103 17 169 93
rect 349 201 431 325
rect 681 441 757 527
rect 975 383 1041 527
rect 1464 451 1540 527
rect 286 17 357 93
rect 717 193 783 213
rect 717 147 799 193
rect 1728 451 2006 527
rect 717 17 751 105
rect 1456 147 1565 213
rect 2040 326 2097 493
rect 1847 219 1938 265
rect 1065 17 1135 93
rect 1450 17 1515 105
rect 1945 17 2006 161
rect 2061 143 2097 326
rect 2040 51 2097 143
rect 2231 353 2289 527
rect 2323 291 2375 493
rect 2333 165 2375 291
rect 2230 17 2289 109
rect 2323 51 2375 165
rect 0 -17 2392 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 168 393
rect 122 187 168 359
rect 35 153 122 161
rect 156 153 168 187
rect 35 127 168 153
rect 203 391 247 493
rect 391 393 425 493
rect 467 450 633 484
rect 203 357 213 391
rect 35 69 69 127
rect 203 69 247 357
rect 281 359 425 393
rect 281 165 315 359
rect 465 357 489 391
rect 523 357 565 391
rect 465 315 565 357
rect 281 127 425 165
rect 465 141 509 315
rect 599 281 633 450
rect 817 407 851 475
rect 667 357 937 407
rect 1250 450 1416 484
rect 1212 391 1259 397
rect 667 315 717 357
rect 819 281 869 297
rect 599 247 869 281
rect 599 239 683 247
rect 545 187 615 203
rect 545 153 581 187
rect 545 129 615 153
rect 391 61 425 127
rect 649 93 683 239
rect 825 231 869 247
rect 903 213 937 357
rect 1212 357 1225 391
rect 971 323 1172 331
rect 971 289 1133 323
rect 1167 289 1172 323
rect 1212 315 1259 357
rect 971 283 1172 289
rect 971 247 1037 283
rect 1307 261 1348 381
rect 1213 255 1348 261
rect 1099 213 1165 247
rect 903 179 1165 213
rect 1213 221 1225 255
rect 1259 225 1348 255
rect 1382 281 1416 450
rect 1588 417 1622 475
rect 1450 383 2006 417
rect 1450 315 1500 383
rect 1382 247 1652 281
rect 1259 221 1281 225
rect 1213 212 1281 221
rect 903 153 947 179
rect 881 119 947 153
rect 480 53 683 93
rect 785 85 851 101
rect 981 85 1015 143
rect 1237 141 1281 212
rect 1382 93 1416 247
rect 1608 215 1652 247
rect 1686 168 1720 383
rect 1754 323 1911 349
rect 1754 289 1771 323
rect 1805 315 1911 323
rect 1805 289 1811 315
rect 1754 222 1811 289
rect 1972 265 2006 383
rect 1767 185 1811 222
rect 1972 199 2025 265
rect 1686 167 1723 168
rect 1643 133 1723 167
rect 1767 151 1895 185
rect 785 51 1015 85
rect 1260 53 1416 93
rect 1549 85 1615 109
rect 1757 85 1791 117
rect 1549 51 1791 85
rect 1853 53 1895 151
rect 2132 265 2195 483
rect 2132 199 2299 265
rect 2132 51 2195 199
<< obsli1c >>
rect 122 153 156 187
rect 213 357 247 391
rect 489 357 523 391
rect 581 153 615 187
rect 1225 357 1259 391
rect 1133 289 1167 323
rect 1225 221 1259 255
rect 1771 289 1805 323
<< metal1 >>
rect 0 496 2392 592
rect 753 184 811 193
rect 1503 184 1561 193
rect 753 156 1561 184
rect 753 147 811 156
rect 1503 147 1561 156
rect 0 -48 2392 48
<< obsm1 >>
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 477 391 535 397
rect 477 388 489 391
rect 247 360 489 388
rect 247 357 259 360
rect 201 351 259 357
rect 477 357 489 360
rect 523 388 535 391
rect 1213 391 1271 397
rect 1213 388 1225 391
rect 523 360 1225 388
rect 523 357 535 360
rect 477 351 535 357
rect 1213 357 1225 360
rect 1259 357 1271 391
rect 1213 351 1271 357
rect 1121 323 1179 329
rect 1121 289 1133 323
rect 1167 320 1179 323
rect 1759 323 1817 329
rect 1759 320 1771 323
rect 1167 292 1771 320
rect 1167 289 1179 292
rect 1121 283 1179 289
rect 1759 289 1771 292
rect 1805 289 1817 323
rect 1759 283 1817 289
rect 1213 255 1271 261
rect 1213 252 1225 255
rect 584 224 1225 252
rect 584 193 627 224
rect 1213 221 1225 224
rect 1259 221 1271 255
rect 1213 215 1271 221
rect 110 187 168 193
rect 110 153 122 187
rect 156 184 168 187
rect 569 187 627 193
rect 569 184 581 187
rect 156 156 581 184
rect 156 153 168 156
rect 110 147 168 153
rect 569 153 581 156
rect 615 153 627 187
rect 569 147 627 153
<< labels >>
rlabel locali s 349 201 431 325 6 D
port 1 nsew signal input
rlabel locali s 2333 165 2375 291 6 Q
port 2 nsew signal output
rlabel locali s 2323 291 2375 493 6 Q
port 2 nsew signal output
rlabel locali s 2323 51 2375 165 6 Q
port 2 nsew signal output
rlabel locali s 2061 143 2097 326 6 Q_N
port 3 nsew signal output
rlabel locali s 2040 326 2097 493 6 Q_N
port 3 nsew signal output
rlabel locali s 2040 51 2097 143 6 Q_N
port 3 nsew signal output
rlabel locali s 1847 219 1938 265 6 RESET_B
port 4 nsew signal input
rlabel locali s 717 193 783 213 6 SET_B
port 5 nsew signal input
rlabel locali s 717 147 799 193 6 SET_B
port 5 nsew signal input
rlabel locali s 1456 147 1565 213 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1503 184 1561 193 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1503 147 1561 156 6 SET_B
port 5 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 5 nsew signal input
rlabel metal1 s 753 156 1561 184 6 SET_B
port 5 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 5 nsew signal input
rlabel locali s 17 195 87 325 6 CLK_N
port 6 nsew clock input
rlabel locali s 2230 17 2289 109 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1945 17 2006 161 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1450 17 1515 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 1065 17 1135 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 717 17 751 105 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 286 17 357 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 2392 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2392 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 2231 353 2289 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1728 451 2006 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1464 451 1540 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 975 383 1041 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 681 441 757 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 286 427 357 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 2392 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 2392 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3319692
string GDS_START 3300142
<< end >>
