magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 17 297 76 527
rect 110 263 181 493
rect 215 367 294 527
rect 17 211 181 263
rect 110 199 181 211
rect 396 265 450 414
rect 283 199 350 265
rect 384 199 450 265
rect 488 265 535 414
rect 672 367 719 527
rect 488 199 546 265
rect 580 199 660 265
rect 17 17 76 177
rect 110 51 165 199
rect 762 199 811 265
rect 199 17 333 165
rect 460 17 535 97
rect 0 -17 828 17
<< obsli1 >>
rect 328 459 635 493
rect 328 333 362 459
rect 215 299 362 333
rect 215 199 249 299
rect 569 333 635 459
rect 753 333 811 493
rect 569 299 811 333
rect 694 165 728 299
rect 367 131 644 165
rect 367 62 424 131
rect 578 62 644 131
rect 694 51 811 165
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 283 199 350 265 6 A1
port 1 nsew signal input
rlabel locali s 396 265 450 414 6 A2
port 2 nsew signal input
rlabel locali s 384 199 450 265 6 A2
port 2 nsew signal input
rlabel locali s 488 265 535 414 6 A3
port 3 nsew signal input
rlabel locali s 488 199 546 265 6 A3
port 3 nsew signal input
rlabel locali s 580 199 660 265 6 B1
port 4 nsew signal input
rlabel locali s 762 199 811 265 6 C1
port 5 nsew signal input
rlabel locali s 110 263 181 493 6 X
port 6 nsew signal output
rlabel locali s 110 199 181 211 6 X
port 6 nsew signal output
rlabel locali s 110 51 165 199 6 X
port 6 nsew signal output
rlabel locali s 17 211 181 263 6 X
port 6 nsew signal output
rlabel locali s 460 17 535 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 199 17 333 165 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 17 17 76 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 672 367 719 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 215 367 294 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 297 76 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 755820
string GDS_START 747470
<< end >>
