magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scnmos >>
rect 99 74 129 222
rect 215 94 245 222
rect 315 94 345 222
rect 529 74 559 202
rect 615 74 645 202
rect 715 74 745 202
<< pmoshvt >>
rect 86 368 116 592
rect 234 392 264 592
rect 318 392 348 592
rect 432 392 462 592
rect 546 392 576 592
rect 748 392 778 592
<< ndiff >>
rect 42 210 99 222
rect 42 176 54 210
rect 88 176 99 210
rect 42 120 99 176
rect 42 86 54 120
rect 88 86 99 120
rect 42 74 99 86
rect 129 210 215 222
rect 129 176 154 210
rect 188 176 215 210
rect 129 120 215 176
rect 129 86 154 120
rect 188 94 215 120
rect 245 210 315 222
rect 245 176 256 210
rect 290 176 315 210
rect 245 140 315 176
rect 245 106 256 140
rect 290 106 315 140
rect 245 94 315 106
rect 345 164 402 222
rect 345 130 356 164
rect 390 130 402 164
rect 345 94 402 130
rect 456 188 529 202
rect 456 154 468 188
rect 502 154 529 188
rect 456 120 529 154
rect 188 86 200 94
rect 129 74 200 86
rect 456 86 484 120
rect 518 86 529 120
rect 456 74 529 86
rect 559 179 615 202
rect 559 145 570 179
rect 604 145 615 179
rect 559 74 615 145
rect 645 190 715 202
rect 645 156 670 190
rect 704 156 715 190
rect 645 122 715 156
rect 645 88 670 122
rect 704 88 715 122
rect 645 74 715 88
rect 745 190 837 202
rect 745 156 770 190
rect 804 156 837 190
rect 745 122 837 156
rect 745 88 770 122
rect 804 88 837 122
rect 745 74 837 88
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 234 592
rect 116 546 157 580
rect 191 546 234 580
rect 116 500 234 546
rect 116 466 157 500
rect 191 466 234 500
rect 116 392 234 466
rect 264 392 318 592
rect 348 580 432 592
rect 348 546 361 580
rect 395 546 432 580
rect 348 510 432 546
rect 348 476 361 510
rect 395 476 432 510
rect 348 440 432 476
rect 348 406 361 440
rect 395 406 432 440
rect 348 392 432 406
rect 462 392 546 592
rect 576 580 748 592
rect 576 546 589 580
rect 623 546 691 580
rect 725 546 748 580
rect 576 494 748 546
rect 576 460 589 494
rect 623 460 691 494
rect 725 460 748 494
rect 576 392 748 460
rect 778 580 837 592
rect 778 546 791 580
rect 825 546 837 580
rect 778 511 837 546
rect 778 477 791 511
rect 825 477 837 511
rect 778 442 837 477
rect 778 408 791 442
rect 825 408 837 442
rect 778 392 837 408
rect 116 368 169 392
<< ndiffc >>
rect 54 176 88 210
rect 54 86 88 120
rect 154 176 188 210
rect 154 86 188 120
rect 256 176 290 210
rect 256 106 290 140
rect 356 130 390 164
rect 468 154 502 188
rect 484 86 518 120
rect 570 145 604 179
rect 670 156 704 190
rect 670 88 704 122
rect 770 156 804 190
rect 770 88 804 122
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 157 546 191 580
rect 157 466 191 500
rect 361 546 395 580
rect 361 476 395 510
rect 361 406 395 440
rect 589 546 623 580
rect 691 546 725 580
rect 589 460 623 494
rect 691 460 725 494
rect 791 546 825 580
rect 791 477 825 511
rect 791 408 825 442
<< poly >>
rect 86 592 116 618
rect 234 592 264 618
rect 318 592 348 618
rect 432 592 462 618
rect 546 592 576 618
rect 748 592 778 618
rect 234 377 264 392
rect 318 377 348 392
rect 432 377 462 392
rect 546 377 576 392
rect 748 377 778 392
rect 86 353 116 368
rect 231 356 267 377
rect 83 330 119 353
rect 201 340 267 356
rect 83 314 157 330
rect 83 280 107 314
rect 141 280 157 314
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 315 356 351 377
rect 429 356 465 377
rect 543 358 579 377
rect 745 358 781 377
rect 315 340 381 356
rect 315 306 331 340
rect 365 306 381 340
rect 315 290 381 306
rect 429 340 495 356
rect 429 306 445 340
rect 479 306 495 340
rect 543 342 651 358
rect 543 328 601 342
rect 83 264 157 280
rect 99 222 129 264
rect 215 222 245 290
rect 315 222 345 290
rect 429 250 495 306
rect 585 308 601 328
rect 635 308 651 342
rect 585 292 651 308
rect 699 342 781 358
rect 699 308 715 342
rect 749 308 781 342
rect 429 220 559 250
rect 529 202 559 220
rect 615 202 645 292
rect 699 274 781 308
rect 699 240 715 274
rect 749 240 781 274
rect 699 224 781 240
rect 715 202 745 224
rect 99 48 129 74
rect 215 68 245 94
rect 315 68 345 94
rect 529 48 559 74
rect 615 48 645 74
rect 715 48 745 74
<< polycont >>
rect 107 280 141 314
rect 217 306 251 340
rect 331 306 365 340
rect 445 306 479 340
rect 601 308 635 342
rect 715 308 749 342
rect 715 240 749 274
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 136 580 212 649
rect 136 546 157 580
rect 191 546 212 580
rect 136 500 212 546
rect 136 466 157 500
rect 191 466 212 500
rect 136 458 212 466
rect 345 580 411 596
rect 345 546 361 580
rect 395 546 411 580
rect 345 510 411 546
rect 345 476 361 510
rect 395 476 411 510
rect 345 440 411 476
rect 573 580 741 649
rect 573 546 589 580
rect 623 546 691 580
rect 725 546 741 580
rect 573 494 741 546
rect 573 460 589 494
rect 623 460 691 494
rect 725 460 741 494
rect 775 580 841 596
rect 775 546 791 580
rect 825 546 841 580
rect 775 511 841 546
rect 775 477 791 511
rect 825 477 841 511
rect 345 424 361 440
rect 23 380 39 414
rect 73 380 89 414
rect 23 364 89 380
rect 123 406 361 424
rect 395 426 411 440
rect 775 442 841 477
rect 775 426 791 442
rect 395 408 791 426
rect 825 408 841 442
rect 395 406 841 408
rect 123 392 841 406
rect 123 390 411 392
rect 23 226 57 364
rect 123 330 157 390
rect 91 314 157 330
rect 91 280 107 314
rect 141 280 157 314
rect 201 340 267 356
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 313 340 381 356
rect 313 306 331 340
rect 365 306 381 340
rect 313 290 381 306
rect 429 340 551 356
rect 429 306 445 340
rect 479 306 551 340
rect 429 290 551 306
rect 585 342 651 358
rect 585 308 601 342
rect 635 308 651 342
rect 585 292 651 308
rect 697 342 765 358
rect 697 308 715 342
rect 749 308 765 342
rect 91 264 157 280
rect 697 274 765 308
rect 23 210 104 226
rect 23 176 54 210
rect 88 176 104 210
rect 23 120 104 176
rect 23 86 54 120
rect 88 86 104 120
rect 23 70 104 86
rect 138 210 204 226
rect 138 176 154 210
rect 188 176 204 210
rect 138 120 204 176
rect 138 86 154 120
rect 188 86 204 120
rect 240 222 620 256
rect 697 240 715 274
rect 749 240 765 274
rect 697 224 765 240
rect 240 210 306 222
rect 240 176 256 210
rect 290 176 306 210
rect 240 140 306 176
rect 240 106 256 140
rect 290 106 306 140
rect 240 90 306 106
rect 340 164 406 188
rect 340 130 356 164
rect 390 130 406 164
rect 138 17 204 86
rect 340 17 406 130
rect 452 154 468 188
rect 502 154 518 188
rect 452 120 518 154
rect 452 86 484 120
rect 554 179 620 222
rect 807 190 841 392
rect 554 145 570 179
rect 604 145 620 179
rect 554 119 620 145
rect 654 156 670 190
rect 704 156 720 190
rect 654 122 720 156
rect 452 85 518 86
rect 654 88 670 122
rect 704 88 720 122
rect 654 85 720 88
rect 452 51 720 85
rect 754 156 770 190
rect 804 156 841 190
rect 754 122 841 156
rect 754 88 770 122
rect 804 88 841 122
rect 754 72 841 88
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o221a_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 864 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1520992
string GDS_START 1513042
<< end >>
