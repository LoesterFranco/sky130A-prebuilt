magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 281 47 311 177
rect 365 47 395 177
rect 459 47 489 177
rect 553 47 583 177
rect 647 47 677 177
rect 741 47 771 177
rect 845 47 875 177
rect 1050 47 1080 177
rect 1144 47 1174 177
rect 1238 47 1268 177
rect 1332 47 1362 177
rect 1426 47 1456 177
rect 1520 47 1550 177
rect 1614 47 1644 177
rect 1708 47 1738 177
<< pmoshvt >>
rect 81 297 117 497
rect 289 309 325 497
rect 383 309 419 497
rect 477 309 513 497
rect 571 309 607 497
rect 665 309 701 497
rect 759 309 795 497
rect 853 309 889 497
rect 947 309 983 497
rect 1052 297 1088 497
rect 1146 297 1182 497
rect 1240 297 1276 497
rect 1334 297 1370 497
rect 1428 297 1464 497
rect 1522 297 1558 497
rect 1616 297 1652 497
rect 1710 297 1746 497
<< ndiff >>
rect 27 106 79 177
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 183 177
rect 109 55 129 89
rect 163 55 183 89
rect 109 47 183 55
rect 213 124 281 177
rect 213 90 227 124
rect 261 90 281 124
rect 213 47 281 90
rect 311 89 365 177
rect 311 55 321 89
rect 355 55 365 89
rect 311 47 365 55
rect 395 124 459 177
rect 395 90 415 124
rect 449 90 459 124
rect 395 47 459 90
rect 489 89 553 177
rect 489 55 509 89
rect 543 55 553 89
rect 489 47 553 55
rect 583 124 647 177
rect 583 90 603 124
rect 637 90 647 124
rect 583 47 647 90
rect 677 89 741 177
rect 677 55 697 89
rect 731 55 741 89
rect 677 47 741 55
rect 771 124 845 177
rect 771 90 791 124
rect 825 90 845 124
rect 771 47 845 90
rect 875 89 931 177
rect 875 55 885 89
rect 919 55 931 89
rect 875 47 931 55
rect 998 124 1050 177
rect 998 90 1006 124
rect 1040 90 1050 124
rect 998 47 1050 90
rect 1080 169 1144 177
rect 1080 135 1100 169
rect 1134 135 1144 169
rect 1080 47 1144 135
rect 1174 89 1238 177
rect 1174 55 1194 89
rect 1228 55 1238 89
rect 1174 47 1238 55
rect 1268 169 1332 177
rect 1268 135 1288 169
rect 1322 135 1332 169
rect 1268 47 1332 135
rect 1362 89 1426 177
rect 1362 55 1382 89
rect 1416 55 1426 89
rect 1362 47 1426 55
rect 1456 169 1520 177
rect 1456 135 1476 169
rect 1510 135 1520 169
rect 1456 47 1520 135
rect 1550 89 1614 177
rect 1550 55 1570 89
rect 1604 55 1614 89
rect 1550 47 1614 55
rect 1644 169 1708 177
rect 1644 135 1664 169
rect 1698 135 1708 169
rect 1644 47 1708 135
rect 1738 89 1804 177
rect 1738 55 1758 89
rect 1792 55 1804 89
rect 1738 47 1804 55
<< pdiff >>
rect 27 450 81 497
rect 27 416 35 450
rect 69 416 81 450
rect 27 297 81 416
rect 117 485 171 497
rect 117 451 129 485
rect 163 451 171 485
rect 117 297 171 451
rect 235 465 289 497
rect 235 431 243 465
rect 277 431 289 465
rect 235 309 289 431
rect 325 489 383 497
rect 325 455 337 489
rect 371 455 383 489
rect 325 421 383 455
rect 325 387 337 421
rect 371 387 383 421
rect 325 309 383 387
rect 419 477 477 497
rect 419 443 431 477
rect 465 443 477 477
rect 419 409 477 443
rect 419 375 431 409
rect 465 375 477 409
rect 419 309 477 375
rect 513 489 571 497
rect 513 455 525 489
rect 559 455 571 489
rect 513 421 571 455
rect 513 387 525 421
rect 559 387 571 421
rect 513 309 571 387
rect 607 477 665 497
rect 607 443 619 477
rect 653 443 665 477
rect 607 409 665 443
rect 607 375 619 409
rect 653 375 665 409
rect 607 309 665 375
rect 701 489 759 497
rect 701 455 713 489
rect 747 455 759 489
rect 701 421 759 455
rect 701 387 713 421
rect 747 387 759 421
rect 701 309 759 387
rect 795 477 853 497
rect 795 443 807 477
rect 841 443 853 477
rect 795 409 853 443
rect 795 375 807 409
rect 841 375 853 409
rect 795 309 853 375
rect 889 489 947 497
rect 889 455 901 489
rect 935 455 947 489
rect 889 421 947 455
rect 889 387 901 421
rect 935 387 947 421
rect 889 309 947 387
rect 983 477 1052 497
rect 983 443 1001 477
rect 1035 443 1052 477
rect 983 409 1052 443
rect 983 375 1001 409
rect 1035 375 1052 409
rect 983 309 1052 375
rect 1000 297 1052 309
rect 1088 407 1146 497
rect 1088 373 1100 407
rect 1134 373 1146 407
rect 1088 339 1146 373
rect 1088 305 1100 339
rect 1134 305 1146 339
rect 1088 297 1146 305
rect 1182 477 1240 497
rect 1182 443 1194 477
rect 1228 443 1240 477
rect 1182 409 1240 443
rect 1182 375 1194 409
rect 1228 375 1240 409
rect 1182 297 1240 375
rect 1276 407 1334 497
rect 1276 373 1288 407
rect 1322 373 1334 407
rect 1276 339 1334 373
rect 1276 305 1288 339
rect 1322 305 1334 339
rect 1276 297 1334 305
rect 1370 477 1428 497
rect 1370 443 1382 477
rect 1416 443 1428 477
rect 1370 409 1428 443
rect 1370 375 1382 409
rect 1416 375 1428 409
rect 1370 297 1428 375
rect 1464 407 1522 497
rect 1464 373 1476 407
rect 1510 373 1522 407
rect 1464 339 1522 373
rect 1464 305 1476 339
rect 1510 305 1522 339
rect 1464 297 1522 305
rect 1558 477 1616 497
rect 1558 443 1570 477
rect 1604 443 1616 477
rect 1558 409 1616 443
rect 1558 375 1570 409
rect 1604 375 1616 409
rect 1558 297 1616 375
rect 1652 407 1710 497
rect 1652 373 1664 407
rect 1698 373 1710 407
rect 1652 339 1710 373
rect 1652 305 1664 339
rect 1698 305 1710 339
rect 1652 297 1710 305
rect 1746 477 1800 497
rect 1746 443 1758 477
rect 1792 443 1800 477
rect 1746 409 1800 443
rect 1746 375 1758 409
rect 1792 375 1800 409
rect 1746 297 1800 375
<< ndiffc >>
rect 35 72 69 106
rect 129 55 163 89
rect 227 90 261 124
rect 321 55 355 89
rect 415 90 449 124
rect 509 55 543 89
rect 603 90 637 124
rect 697 55 731 89
rect 791 90 825 124
rect 885 55 919 89
rect 1006 90 1040 124
rect 1100 135 1134 169
rect 1194 55 1228 89
rect 1288 135 1322 169
rect 1382 55 1416 89
rect 1476 135 1510 169
rect 1570 55 1604 89
rect 1664 135 1698 169
rect 1758 55 1792 89
<< pdiffc >>
rect 35 416 69 450
rect 129 451 163 485
rect 243 431 277 465
rect 337 455 371 489
rect 337 387 371 421
rect 431 443 465 477
rect 431 375 465 409
rect 525 455 559 489
rect 525 387 559 421
rect 619 443 653 477
rect 619 375 653 409
rect 713 455 747 489
rect 713 387 747 421
rect 807 443 841 477
rect 807 375 841 409
rect 901 455 935 489
rect 901 387 935 421
rect 1001 443 1035 477
rect 1001 375 1035 409
rect 1100 373 1134 407
rect 1100 305 1134 339
rect 1194 443 1228 477
rect 1194 375 1228 409
rect 1288 373 1322 407
rect 1288 305 1322 339
rect 1382 443 1416 477
rect 1382 375 1416 409
rect 1476 373 1510 407
rect 1476 305 1510 339
rect 1570 443 1604 477
rect 1570 375 1604 409
rect 1664 373 1698 407
rect 1664 305 1698 339
rect 1758 443 1792 477
rect 1758 375 1792 409
<< poly >>
rect 81 497 117 523
rect 289 497 325 523
rect 383 497 419 523
rect 477 497 513 523
rect 571 497 607 523
rect 665 497 701 523
rect 759 497 795 523
rect 853 497 889 523
rect 947 497 983 523
rect 1052 497 1088 523
rect 1146 497 1182 523
rect 1240 497 1276 523
rect 1334 497 1370 523
rect 1428 497 1464 523
rect 1522 497 1558 523
rect 1616 497 1652 523
rect 1710 497 1746 523
rect 81 282 117 297
rect 289 294 325 309
rect 383 294 419 309
rect 477 294 513 309
rect 571 294 607 309
rect 665 294 701 309
rect 759 294 795 309
rect 853 294 889 309
rect 947 294 983 309
rect 79 265 119 282
rect 22 249 119 265
rect 287 264 985 294
rect 1052 282 1088 297
rect 1146 282 1182 297
rect 1240 282 1276 297
rect 1334 282 1370 297
rect 1428 282 1464 297
rect 1522 282 1558 297
rect 1616 282 1652 297
rect 1710 282 1746 297
rect 22 215 32 249
rect 66 222 119 249
rect 921 249 985 264
rect 66 215 875 222
rect 22 199 875 215
rect 921 215 931 249
rect 965 215 985 249
rect 921 199 985 215
rect 1050 265 1090 282
rect 1144 265 1184 282
rect 1050 259 1184 265
rect 1238 259 1278 282
rect 1332 259 1372 282
rect 1426 265 1466 282
rect 1520 265 1560 282
rect 1426 259 1560 265
rect 1614 259 1654 282
rect 1708 261 1748 282
rect 1708 259 1806 261
rect 1050 249 1806 259
rect 1050 215 1220 249
rect 1254 215 1298 249
rect 1332 215 1376 249
rect 1410 215 1444 249
rect 1478 215 1522 249
rect 1556 215 1600 249
rect 1634 215 1678 249
rect 1712 215 1756 249
rect 1790 215 1806 249
rect 1050 205 1806 215
rect 1050 199 1174 205
rect 79 192 875 199
rect 79 177 109 192
rect 183 177 213 192
rect 281 177 311 192
rect 365 177 395 192
rect 459 177 489 192
rect 553 177 583 192
rect 647 177 677 192
rect 741 177 771 192
rect 845 177 875 192
rect 1050 177 1080 199
rect 1144 177 1174 199
rect 1238 177 1268 205
rect 1332 177 1362 205
rect 1426 199 1550 205
rect 1426 177 1456 199
rect 1520 177 1550 199
rect 1614 177 1644 205
rect 1708 203 1806 205
rect 1708 177 1738 203
rect 79 21 109 47
rect 183 21 213 47
rect 281 21 311 47
rect 365 21 395 47
rect 459 21 489 47
rect 553 21 583 47
rect 647 21 677 47
rect 741 21 771 47
rect 845 21 875 47
rect 1050 21 1080 47
rect 1144 21 1174 47
rect 1238 21 1268 47
rect 1332 21 1362 47
rect 1426 21 1456 47
rect 1520 21 1550 47
rect 1614 21 1644 47
rect 1708 21 1738 47
<< polycont >>
rect 32 215 66 249
rect 931 215 965 249
rect 1220 215 1254 249
rect 1298 215 1332 249
rect 1376 215 1410 249
rect 1444 215 1478 249
rect 1522 215 1556 249
rect 1600 215 1634 249
rect 1678 215 1712 249
rect 1756 215 1790 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 17 450 69 493
rect 17 416 35 450
rect 103 485 185 527
rect 103 451 129 485
rect 163 451 185 485
rect 103 425 185 451
rect 235 465 277 493
rect 235 431 243 465
rect 17 391 69 416
rect 17 357 185 391
rect 17 249 66 323
rect 17 215 32 249
rect 17 199 66 215
rect 100 265 185 357
rect 235 345 277 431
rect 321 489 387 527
rect 321 455 337 489
rect 371 455 387 489
rect 321 421 387 455
rect 321 387 337 421
rect 371 387 387 421
rect 321 379 387 387
rect 431 477 465 493
rect 431 409 465 443
rect 509 489 575 527
rect 509 455 525 489
rect 559 455 575 489
rect 509 421 575 455
rect 509 387 525 421
rect 559 387 575 421
rect 509 379 575 387
rect 619 477 653 493
rect 619 409 653 443
rect 431 345 465 375
rect 697 489 763 527
rect 697 455 713 489
rect 747 455 763 489
rect 697 421 763 455
rect 697 387 713 421
rect 747 387 763 421
rect 697 379 763 387
rect 807 477 841 493
rect 807 409 841 443
rect 619 345 653 375
rect 885 489 951 527
rect 885 455 901 489
rect 935 455 951 489
rect 885 421 951 455
rect 885 387 901 421
rect 935 387 951 421
rect 885 379 951 387
rect 995 477 1819 493
rect 995 443 1001 477
rect 1035 459 1194 477
rect 1035 443 1040 459
rect 995 409 1040 443
rect 1228 459 1382 477
rect 807 345 841 375
rect 995 375 1001 409
rect 1035 375 1040 409
rect 995 345 1040 375
rect 235 311 1040 345
rect 1074 407 1150 425
rect 1074 373 1100 407
rect 1134 373 1150 407
rect 1074 339 1150 373
rect 1194 409 1228 443
rect 1416 459 1570 477
rect 1194 357 1228 375
rect 1262 407 1338 425
rect 1262 373 1288 407
rect 1322 373 1338 407
rect 1074 305 1100 339
rect 1134 323 1150 339
rect 1262 339 1338 373
rect 1382 409 1416 443
rect 1604 459 1758 477
rect 1382 357 1416 375
rect 1450 407 1526 425
rect 1450 373 1476 407
rect 1510 373 1526 407
rect 1262 323 1288 339
rect 1134 305 1288 323
rect 1322 323 1338 339
rect 1450 339 1526 373
rect 1570 409 1604 443
rect 1792 443 1819 477
rect 1570 357 1604 375
rect 1638 407 1714 425
rect 1638 373 1664 407
rect 1698 373 1714 407
rect 1450 323 1476 339
rect 1322 305 1476 323
rect 1510 323 1526 339
rect 1638 339 1714 373
rect 1638 323 1664 339
rect 1510 305 1664 323
rect 1698 305 1714 339
rect 1074 289 1714 305
rect 1758 409 1819 443
rect 1792 375 1819 409
rect 1758 289 1819 375
rect 100 249 1040 265
rect 100 215 931 249
rect 965 215 1040 249
rect 100 199 1040 215
rect 100 165 149 199
rect 1074 170 1160 289
rect 1204 249 1810 255
rect 1204 215 1220 249
rect 1254 215 1298 249
rect 1332 215 1376 249
rect 1410 215 1444 249
rect 1478 215 1522 249
rect 1556 215 1600 249
rect 1634 215 1678 249
rect 1712 215 1756 249
rect 1790 215 1810 249
rect 1204 204 1810 215
rect 1074 169 1819 170
rect 17 131 149 165
rect 227 131 1040 165
rect 17 106 69 131
rect 17 72 35 106
rect 227 124 261 131
rect 17 51 69 72
rect 103 89 179 97
rect 103 55 129 89
rect 163 55 179 89
rect 103 17 179 55
rect 415 124 449 131
rect 227 51 261 90
rect 295 89 371 97
rect 295 55 321 89
rect 355 55 371 89
rect 295 17 371 55
rect 603 124 637 131
rect 415 51 449 90
rect 483 89 559 97
rect 483 55 509 89
rect 543 55 559 89
rect 483 17 559 55
rect 791 124 825 131
rect 603 51 637 90
rect 671 89 747 97
rect 671 55 697 89
rect 731 55 747 89
rect 671 17 747 55
rect 971 124 1040 131
rect 1074 135 1100 169
rect 1134 135 1288 169
rect 1322 135 1476 169
rect 1510 135 1664 169
rect 1698 135 1819 169
rect 1074 127 1819 135
rect 791 51 825 90
rect 859 89 937 97
rect 859 55 885 89
rect 919 55 937 89
rect 859 17 937 55
rect 971 90 1006 124
rect 1040 90 1819 93
rect 971 89 1819 90
rect 971 55 1194 89
rect 1228 55 1382 89
rect 1416 55 1570 89
rect 1604 55 1758 89
rect 1792 55 1819 89
rect 971 51 1819 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1226 221 1260 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1595 221 1629 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1504 221 1538 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1407 221 1441 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1676 289 1710 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1489 357 1523 391 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1523 306 1523 306 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1410 289 1444 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 TE
port 2 nsew
flabel corelocali s 30 289 64 323 0 FreeSans 200 0 0 0 TE
port 2 nsew
flabel corelocali s 1133 289 1167 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1316 289 1350 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1226 289 1260 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1683 221 1717 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1768 221 1802 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 1676 357 1710 391 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel corelocali s 1580 289 1614 323 0 FreeSans 200 0 0 0 Z
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2071196
string GDS_START 2057916
<< end >>
