magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 92 53 122 137
rect 186 53 216 137
rect 280 53 310 137
rect 416 47 446 177
rect 520 47 550 177
<< pmoshvt >>
rect 84 297 120 381
rect 166 297 202 381
rect 272 297 308 381
rect 418 297 454 497
rect 512 297 548 497
<< ndiff >>
rect 325 137 416 177
rect 30 111 92 137
rect 30 77 38 111
rect 72 77 92 111
rect 30 53 92 77
rect 122 97 186 137
rect 122 63 132 97
rect 166 63 186 97
rect 122 53 186 63
rect 216 111 280 137
rect 216 77 226 111
rect 260 77 280 111
rect 216 53 280 77
rect 310 97 416 137
rect 310 63 330 97
rect 364 63 416 97
rect 310 53 416 63
rect 325 47 416 53
rect 446 135 520 177
rect 446 101 466 135
rect 500 101 520 135
rect 446 47 520 101
rect 550 165 607 177
rect 550 131 565 165
rect 599 131 607 165
rect 550 97 607 131
rect 550 63 565 97
rect 599 63 607 97
rect 550 47 607 63
<< pdiff >>
rect 325 485 418 497
rect 325 451 333 485
rect 367 451 418 485
rect 325 417 418 451
rect 325 383 333 417
rect 367 383 418 417
rect 325 381 418 383
rect 30 354 84 381
rect 30 320 38 354
rect 72 320 84 354
rect 30 297 84 320
rect 120 297 166 381
rect 202 297 272 381
rect 308 297 418 381
rect 454 454 512 497
rect 454 420 466 454
rect 500 420 512 454
rect 454 386 512 420
rect 454 352 466 386
rect 500 352 512 386
rect 454 297 512 352
rect 548 477 613 497
rect 548 443 565 477
rect 599 443 613 477
rect 548 409 613 443
rect 548 375 565 409
rect 599 375 613 409
rect 548 341 613 375
rect 548 307 565 341
rect 599 307 613 341
rect 548 297 613 307
<< ndiffc >>
rect 38 77 72 111
rect 132 63 166 97
rect 226 77 260 111
rect 330 63 364 97
rect 466 101 500 135
rect 565 131 599 165
rect 565 63 599 97
<< pdiffc >>
rect 333 451 367 485
rect 333 383 367 417
rect 38 320 72 354
rect 466 420 500 454
rect 466 352 500 386
rect 565 443 599 477
rect 565 375 599 409
rect 565 307 599 341
<< poly >>
rect 418 497 454 523
rect 512 497 548 523
rect 164 473 234 483
rect 164 439 180 473
rect 214 439 234 473
rect 164 429 234 439
rect 164 407 204 429
rect 84 381 120 407
rect 166 381 202 407
rect 272 381 308 407
rect 84 282 120 297
rect 166 282 202 297
rect 272 282 308 297
rect 418 282 454 297
rect 512 282 548 297
rect 82 265 122 282
rect 24 249 122 265
rect 24 215 34 249
rect 68 215 122 249
rect 24 199 122 215
rect 92 137 122 199
rect 164 182 204 282
rect 270 265 310 282
rect 416 265 456 282
rect 510 265 550 282
rect 255 249 319 265
rect 255 215 265 249
rect 299 215 319 249
rect 255 199 319 215
rect 416 249 550 265
rect 416 215 426 249
rect 460 215 550 249
rect 416 199 550 215
rect 164 152 216 182
rect 186 137 216 152
rect 280 137 310 199
rect 416 177 446 199
rect 520 177 550 199
rect 92 27 122 53
rect 186 27 216 53
rect 280 27 310 53
rect 416 21 446 47
rect 520 21 550 47
<< polycont >>
rect 180 439 214 473
rect 34 215 68 249
rect 265 215 299 249
rect 426 215 460 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 320 485 414 527
rect 17 473 276 483
rect 17 439 180 473
rect 214 439 276 473
rect 17 425 276 439
rect 320 451 333 485
rect 367 451 414 485
rect 320 417 414 451
rect 21 357 274 391
rect 320 383 333 417
rect 367 383 414 417
rect 320 367 414 383
rect 466 454 531 493
rect 500 420 531 454
rect 466 386 531 420
rect 21 354 77 357
rect 21 320 38 354
rect 72 320 77 354
rect 240 333 274 357
rect 500 352 531 386
rect 21 299 77 320
rect 111 265 176 323
rect 240 299 422 333
rect 466 299 531 352
rect 378 265 422 299
rect 17 249 77 265
rect 17 215 34 249
rect 68 215 77 249
rect 17 199 77 215
rect 111 249 316 265
rect 111 215 265 249
rect 299 215 316 249
rect 111 199 316 215
rect 378 249 460 265
rect 378 215 426 249
rect 378 199 460 215
rect 378 165 422 199
rect 21 131 422 165
rect 494 152 531 299
rect 565 477 623 527
rect 599 443 623 477
rect 565 409 623 443
rect 599 375 623 409
rect 565 341 623 375
rect 599 307 623 341
rect 565 286 623 307
rect 466 135 531 152
rect 21 111 72 131
rect 21 77 38 111
rect 226 111 260 131
rect 21 61 72 77
rect 106 63 132 97
rect 166 63 182 97
rect 106 17 182 63
rect 500 101 531 135
rect 226 61 260 77
rect 294 63 330 97
rect 364 63 418 97
rect 466 83 531 101
rect 565 165 623 183
rect 599 131 623 165
rect 565 97 623 131
rect 294 17 418 63
rect 599 63 623 97
rect 565 17 623 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel corelocali s 131 221 165 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 216 221 250 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 29 431 63 465 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 475 357 509 391 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel corelocali s 131 289 165 323 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 126 430 160 464 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 217 430 251 464 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 or3_2
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 465000
string GDS_START 458956
<< end >>
