magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 116 367 167 527
rect 207 401 273 493
rect 307 435 422 527
rect 456 401 527 493
rect 207 367 527 401
rect 91 199 160 265
rect 306 181 362 367
rect 398 255 436 331
rect 472 299 527 367
rect 561 299 627 527
rect 398 215 627 255
rect 103 17 169 165
rect 306 161 371 181
rect 305 127 371 161
rect 489 17 523 105
rect 0 -17 644 17
<< obsli1 >>
rect 22 333 82 372
rect 22 299 272 333
rect 22 168 56 299
rect 206 215 272 299
rect 22 102 69 168
rect 216 93 271 181
rect 405 139 627 181
rect 405 93 455 139
rect 216 51 455 93
rect 557 51 627 139
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 91 199 160 265 6 A_N
port 1 nsew signal input
rlabel locali s 398 255 436 331 6 B
port 2 nsew signal input
rlabel locali s 398 215 627 255 6 B
port 2 nsew signal input
rlabel locali s 472 299 527 367 6 Y
port 3 nsew signal output
rlabel locali s 456 401 527 493 6 Y
port 3 nsew signal output
rlabel locali s 306 181 362 367 6 Y
port 3 nsew signal output
rlabel locali s 306 161 371 181 6 Y
port 3 nsew signal output
rlabel locali s 305 127 371 161 6 Y
port 3 nsew signal output
rlabel locali s 207 401 273 493 6 Y
port 3 nsew signal output
rlabel locali s 207 367 527 401 6 Y
port 3 nsew signal output
rlabel locali s 489 17 523 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 165 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 561 299 627 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 307 435 422 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 116 367 167 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1722000
string GDS_START 1715438
<< end >>
