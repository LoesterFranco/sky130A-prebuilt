magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 25 290 110 356
rect 212 290 278 356
rect 586 294 652 360
rect 796 269 873 356
rect 975 394 1041 596
rect 1171 394 1221 596
rect 975 360 1221 394
rect 1171 330 1221 360
rect 1171 296 1319 330
rect 1273 226 1319 296
rect 966 192 1319 226
rect 966 70 1016 192
rect 1152 70 1218 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 390 79 649
rect 203 482 269 649
rect 312 448 346 596
rect 113 390 346 448
rect 144 251 178 390
rect 312 354 346 390
rect 386 388 452 649
rect 486 428 552 596
rect 586 462 729 649
rect 763 428 829 596
rect 863 458 929 649
rect 486 424 829 428
rect 486 394 941 424
rect 486 354 552 394
rect 763 390 941 394
rect 312 320 552 354
rect 907 326 941 390
rect 1081 428 1131 649
rect 1255 364 1321 649
rect 907 260 1137 326
rect 28 97 78 251
rect 144 201 266 251
rect 388 235 762 260
rect 388 226 814 235
rect 114 131 352 167
rect 388 97 422 226
rect 728 199 814 226
rect 458 165 694 192
rect 458 158 728 165
rect 458 115 524 158
rect 28 63 422 97
rect 560 17 626 124
rect 660 115 728 158
rect 866 17 932 226
rect 1052 17 1118 158
rect 1252 17 1304 136
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel locali s 212 290 278 356 6 A
port 1 nsew signal input
rlabel locali s 25 290 110 356 6 B
port 2 nsew signal input
rlabel locali s 796 269 873 356 6 C
port 3 nsew signal input
rlabel locali s 586 294 652 360 6 D
port 4 nsew signal input
rlabel locali s 1273 226 1319 296 6 X
port 5 nsew signal output
rlabel locali s 1171 394 1221 596 6 X
port 5 nsew signal output
rlabel locali s 1171 330 1221 360 6 X
port 5 nsew signal output
rlabel locali s 1171 296 1319 330 6 X
port 5 nsew signal output
rlabel locali s 1152 70 1218 192 6 X
port 5 nsew signal output
rlabel locali s 975 394 1041 596 6 X
port 5 nsew signal output
rlabel locali s 975 360 1221 394 6 X
port 5 nsew signal output
rlabel locali s 966 192 1319 226 6 X
port 5 nsew signal output
rlabel locali s 966 70 1016 192 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1344 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1344 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3213694
string GDS_START 3202796
<< end >>
