magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 356 1670 704
rect -38 332 620 356
rect 979 332 1670 356
<< pwell >>
rect 0 0 1632 49
<< scnmos >>
rect 84 90 114 238
rect 173 90 203 238
rect 289 90 319 238
rect 375 90 405 238
rect 557 110 587 238
rect 643 110 673 238
rect 745 139 775 267
rect 831 139 861 267
rect 1049 122 1079 250
rect 1135 122 1165 250
rect 1221 122 1251 250
rect 1323 122 1353 250
rect 1413 122 1443 250
rect 1518 122 1548 250
<< pmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 276 368 306 592
rect 366 368 396 592
rect 568 392 598 592
rect 668 392 698 592
rect 768 392 798 592
rect 868 392 898 592
rect 1007 392 1037 592
rect 1130 392 1160 592
rect 1224 392 1254 592
rect 1326 392 1356 592
rect 1416 392 1446 592
rect 1516 392 1546 592
<< ndiff >>
rect 688 253 745 267
rect 688 238 700 253
rect 27 136 84 238
rect 27 102 39 136
rect 73 102 84 136
rect 27 90 84 102
rect 114 230 173 238
rect 114 196 126 230
rect 160 196 173 230
rect 114 132 173 196
rect 114 98 126 132
rect 160 98 173 132
rect 114 90 173 98
rect 203 136 289 238
rect 203 102 222 136
rect 256 102 289 136
rect 203 90 289 102
rect 319 220 375 238
rect 319 186 330 220
rect 364 186 375 220
rect 319 136 375 186
rect 319 102 330 136
rect 364 102 375 136
rect 319 90 375 102
rect 405 230 557 238
rect 405 196 430 230
rect 464 196 557 230
rect 405 152 557 196
rect 405 118 430 152
rect 464 118 557 152
rect 405 110 557 118
rect 587 226 643 238
rect 587 192 598 226
rect 632 192 643 226
rect 587 158 643 192
rect 587 124 598 158
rect 632 124 643 158
rect 587 110 643 124
rect 673 219 700 238
rect 734 219 745 253
rect 673 139 745 219
rect 775 185 831 267
rect 775 151 786 185
rect 820 151 831 185
rect 775 139 831 151
rect 861 200 911 267
rect 861 186 932 200
rect 861 152 886 186
rect 920 152 932 186
rect 861 139 932 152
rect 673 110 723 139
rect 992 170 1049 250
rect 992 136 1004 170
rect 1038 136 1049 170
rect 992 122 1049 136
rect 1079 170 1135 250
rect 1079 136 1090 170
rect 1124 136 1135 170
rect 1079 122 1135 136
rect 1165 237 1221 250
rect 1165 203 1176 237
rect 1210 203 1221 237
rect 1165 122 1221 203
rect 1251 238 1323 250
rect 1251 204 1262 238
rect 1296 204 1323 238
rect 1251 169 1323 204
rect 1251 135 1262 169
rect 1296 135 1323 169
rect 1251 122 1323 135
rect 1353 238 1413 250
rect 1353 204 1364 238
rect 1398 204 1413 238
rect 1353 168 1413 204
rect 1353 134 1364 168
rect 1398 134 1413 168
rect 1353 122 1413 134
rect 1443 168 1518 250
rect 1443 134 1456 168
rect 1490 134 1518 168
rect 1443 122 1518 134
rect 1548 238 1605 250
rect 1548 204 1559 238
rect 1593 204 1605 238
rect 1548 168 1605 204
rect 1548 134 1559 168
rect 1593 134 1605 168
rect 1548 122 1605 134
rect 405 90 455 110
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 497 176 546
rect 116 463 129 497
rect 163 463 176 497
rect 116 414 176 463
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 580 276 592
rect 206 546 219 580
rect 253 546 276 580
rect 206 476 276 546
rect 206 442 219 476
rect 253 442 276 476
rect 206 368 276 442
rect 306 584 366 592
rect 306 550 319 584
rect 353 550 366 584
rect 306 498 366 550
rect 306 464 319 498
rect 353 464 366 498
rect 306 420 366 464
rect 306 386 319 420
rect 353 386 366 420
rect 306 368 366 386
rect 396 580 455 592
rect 396 546 409 580
rect 443 546 455 580
rect 396 498 455 546
rect 396 464 409 498
rect 443 464 455 498
rect 396 368 455 464
rect 509 580 568 592
rect 509 546 521 580
rect 555 546 568 580
rect 509 498 568 546
rect 509 464 521 498
rect 555 464 568 498
rect 509 392 568 464
rect 598 538 668 592
rect 598 504 621 538
rect 655 504 668 538
rect 598 440 668 504
rect 598 406 621 440
rect 655 406 668 440
rect 598 392 668 406
rect 698 580 768 592
rect 698 546 721 580
rect 755 546 768 580
rect 698 498 768 546
rect 698 464 721 498
rect 755 464 768 498
rect 698 392 768 464
rect 798 539 868 592
rect 798 505 821 539
rect 855 505 868 539
rect 798 440 868 505
rect 798 406 821 440
rect 855 406 868 440
rect 798 392 868 406
rect 898 580 1007 592
rect 898 546 935 580
rect 969 546 1007 580
rect 898 504 1007 546
rect 898 470 935 504
rect 969 470 1007 504
rect 898 434 1007 470
rect 898 400 935 434
rect 969 400 1007 434
rect 898 392 1007 400
rect 1037 568 1130 592
rect 1037 534 1061 568
rect 1095 534 1130 568
rect 1037 392 1130 534
rect 1160 580 1224 592
rect 1160 546 1173 580
rect 1207 546 1224 580
rect 1160 492 1224 546
rect 1160 458 1173 492
rect 1207 458 1224 492
rect 1160 392 1224 458
rect 1254 576 1326 592
rect 1254 542 1276 576
rect 1310 542 1326 576
rect 1254 392 1326 542
rect 1356 584 1416 592
rect 1356 550 1369 584
rect 1403 550 1416 584
rect 1356 510 1416 550
rect 1356 476 1369 510
rect 1403 476 1416 510
rect 1356 434 1416 476
rect 1356 400 1369 434
rect 1403 400 1416 434
rect 1356 392 1416 400
rect 1446 584 1516 592
rect 1446 550 1459 584
rect 1493 550 1516 584
rect 1446 508 1516 550
rect 1446 474 1459 508
rect 1493 474 1516 508
rect 1446 392 1516 474
rect 1546 580 1605 592
rect 1546 546 1559 580
rect 1593 546 1605 580
rect 1546 510 1605 546
rect 1546 476 1559 510
rect 1593 476 1605 510
rect 1546 440 1605 476
rect 1546 406 1559 440
rect 1593 406 1605 440
rect 1546 392 1605 406
<< ndiffc >>
rect 39 102 73 136
rect 126 196 160 230
rect 126 98 160 132
rect 222 102 256 136
rect 330 186 364 220
rect 330 102 364 136
rect 430 196 464 230
rect 430 118 464 152
rect 598 192 632 226
rect 598 124 632 158
rect 700 219 734 253
rect 786 151 820 185
rect 886 152 920 186
rect 1004 136 1038 170
rect 1090 136 1124 170
rect 1176 203 1210 237
rect 1262 204 1296 238
rect 1262 135 1296 169
rect 1364 204 1398 238
rect 1364 134 1398 168
rect 1456 134 1490 168
rect 1559 204 1593 238
rect 1559 134 1593 168
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 546 253 580
rect 219 442 253 476
rect 319 550 353 584
rect 319 464 353 498
rect 319 386 353 420
rect 409 546 443 580
rect 409 464 443 498
rect 521 546 555 580
rect 521 464 555 498
rect 621 504 655 538
rect 621 406 655 440
rect 721 546 755 580
rect 721 464 755 498
rect 821 505 855 539
rect 821 406 855 440
rect 935 546 969 580
rect 935 470 969 504
rect 935 400 969 434
rect 1061 534 1095 568
rect 1173 546 1207 580
rect 1173 458 1207 492
rect 1276 542 1310 576
rect 1369 550 1403 584
rect 1369 476 1403 510
rect 1369 400 1403 434
rect 1459 550 1493 584
rect 1459 474 1493 508
rect 1559 546 1593 580
rect 1559 476 1593 510
rect 1559 406 1593 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 276 592 306 618
rect 366 592 396 618
rect 568 592 598 618
rect 668 592 698 618
rect 768 592 798 618
rect 868 592 898 618
rect 1007 592 1037 618
rect 1130 592 1160 618
rect 1224 592 1254 618
rect 1326 592 1356 618
rect 1416 592 1446 618
rect 1516 592 1546 618
rect 568 377 598 392
rect 668 377 698 392
rect 768 377 798 392
rect 868 377 898 392
rect 1007 377 1037 392
rect 1130 377 1160 392
rect 1224 377 1254 392
rect 1326 377 1356 392
rect 1416 377 1446 392
rect 1516 377 1546 392
rect 86 353 116 368
rect 176 353 206 368
rect 276 353 306 368
rect 366 353 396 368
rect 565 356 601 377
rect 83 336 119 353
rect 173 336 209 353
rect 273 336 309 353
rect 363 336 399 353
rect 83 320 399 336
rect 83 286 213 320
rect 247 286 281 320
rect 315 286 349 320
rect 383 300 399 320
rect 501 340 601 356
rect 501 306 517 340
rect 551 306 601 340
rect 665 371 701 377
rect 765 371 801 377
rect 665 341 801 371
rect 865 371 901 377
rect 865 341 956 371
rect 665 340 775 341
rect 665 320 681 340
rect 383 286 405 300
rect 501 290 601 306
rect 643 306 681 320
rect 715 306 775 340
rect 643 290 775 306
rect 83 283 405 286
rect 84 270 405 283
rect 84 253 203 270
rect 84 238 114 253
rect 173 238 203 253
rect 289 238 319 270
rect 375 238 405 270
rect 557 238 587 290
rect 643 238 673 290
rect 745 267 775 290
rect 831 267 861 293
rect 926 246 956 341
rect 1004 360 1040 377
rect 1004 344 1079 360
rect 1004 310 1020 344
rect 1054 310 1079 344
rect 1004 294 1079 310
rect 1049 250 1079 294
rect 1127 356 1163 377
rect 1221 356 1257 377
rect 1127 340 1257 356
rect 1323 354 1359 377
rect 1413 356 1449 377
rect 1513 356 1549 377
rect 1127 306 1143 340
rect 1177 306 1257 340
rect 1127 290 1257 306
rect 1299 338 1365 354
rect 1299 304 1315 338
rect 1349 304 1365 338
rect 1135 250 1165 290
rect 1221 250 1251 290
rect 1299 288 1365 304
rect 1413 340 1563 356
rect 1413 306 1429 340
rect 1463 306 1513 340
rect 1547 306 1563 340
rect 1413 290 1563 306
rect 1323 250 1353 288
rect 1413 250 1443 290
rect 1518 250 1548 290
rect 926 216 977 246
rect 745 113 775 139
rect 831 117 861 139
rect 947 117 977 216
rect 84 64 114 90
rect 173 64 203 90
rect 289 64 319 90
rect 375 64 405 90
rect 557 84 587 110
rect 643 84 673 110
rect 817 101 977 117
rect 817 67 833 101
rect 867 87 977 101
rect 1049 96 1079 122
rect 1135 96 1165 122
rect 1221 96 1251 122
rect 1323 96 1353 122
rect 1413 96 1443 122
rect 1518 96 1548 122
rect 867 67 883 87
rect 817 51 883 67
<< polycont >>
rect 213 286 247 320
rect 281 286 315 320
rect 349 286 383 320
rect 517 306 551 340
rect 681 306 715 340
rect 1020 310 1054 344
rect 1143 306 1177 340
rect 1315 304 1349 338
rect 1429 306 1463 340
rect 1513 306 1547 340
rect 833 67 867 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 163 596
rect 113 546 129 580
rect 113 497 163 546
rect 113 463 129 497
rect 113 414 163 463
rect 203 580 269 649
rect 203 546 219 580
rect 253 546 269 580
rect 203 476 269 546
rect 203 442 219 476
rect 253 442 269 476
rect 203 438 269 442
rect 303 584 359 600
rect 303 550 319 584
rect 353 550 359 584
rect 303 498 359 550
rect 303 464 319 498
rect 353 464 359 498
rect 113 380 129 414
rect 303 420 359 464
rect 393 580 459 649
rect 393 546 409 580
rect 443 546 459 580
rect 393 498 459 546
rect 393 464 409 498
rect 443 464 459 498
rect 393 458 459 464
rect 505 581 985 615
rect 505 580 571 581
rect 505 546 521 580
rect 555 546 571 580
rect 705 580 771 581
rect 505 498 571 546
rect 505 464 521 498
rect 555 464 571 498
rect 505 458 571 464
rect 605 538 671 547
rect 605 504 621 538
rect 655 504 671 538
rect 605 440 671 504
rect 705 546 721 580
rect 755 546 771 580
rect 919 580 985 581
rect 705 498 771 546
rect 705 464 721 498
rect 755 464 771 498
rect 705 458 771 464
rect 805 539 871 547
rect 805 505 821 539
rect 855 505 871 539
rect 605 424 621 440
rect 303 404 319 420
rect 163 386 319 404
rect 353 386 359 420
rect 163 380 359 386
rect 113 370 359 380
rect 403 406 621 424
rect 655 424 671 440
rect 805 440 871 505
rect 805 424 821 440
rect 655 406 821 424
rect 855 406 871 440
rect 403 390 871 406
rect 919 546 935 580
rect 969 546 985 580
rect 919 504 985 546
rect 1042 568 1123 649
rect 1042 534 1061 568
rect 1095 534 1123 568
rect 1042 526 1123 534
rect 1157 546 1173 580
rect 1207 546 1223 580
rect 919 470 935 504
rect 969 492 985 504
rect 1157 492 1223 546
rect 1257 576 1329 649
rect 1257 542 1276 576
rect 1310 542 1329 576
rect 1257 526 1329 542
rect 1363 584 1419 600
rect 1363 550 1369 584
rect 1403 550 1419 584
rect 1363 510 1419 550
rect 1363 492 1369 510
rect 969 470 1173 492
rect 919 458 1173 470
rect 1207 476 1369 492
rect 1403 476 1419 510
rect 1207 458 1419 476
rect 1453 584 1509 649
rect 1453 550 1459 584
rect 1493 550 1509 584
rect 1453 508 1509 550
rect 1453 474 1459 508
rect 1493 474 1509 508
rect 1453 458 1509 474
rect 1543 580 1609 596
rect 1543 546 1559 580
rect 1593 546 1609 580
rect 1543 510 1609 546
rect 1543 476 1559 510
rect 1593 476 1609 510
rect 919 434 985 458
rect 919 400 935 434
rect 969 400 985 434
rect 1353 434 1419 458
rect 919 392 985 400
rect 1036 390 1319 424
rect 1353 400 1369 434
rect 1403 424 1419 434
rect 1543 440 1609 476
rect 1543 424 1559 440
rect 1403 406 1559 424
rect 1593 406 1609 440
rect 1403 400 1609 406
rect 1353 390 1609 400
rect 113 330 163 370
rect 403 336 437 390
rect 25 296 163 330
rect 197 320 437 336
rect 25 236 71 296
rect 197 286 213 320
rect 247 286 281 320
rect 315 286 349 320
rect 383 286 437 320
rect 501 340 567 356
rect 501 306 517 340
rect 551 306 567 340
rect 501 290 567 306
rect 601 340 743 356
rect 601 306 681 340
rect 715 306 743 340
rect 601 290 743 306
rect 197 270 437 286
rect 25 230 380 236
rect 25 196 126 230
rect 160 220 380 230
rect 160 196 330 220
rect 25 186 330 196
rect 364 186 380 220
rect 23 136 89 152
rect 23 102 39 136
rect 73 102 89 136
rect 23 17 89 102
rect 123 132 164 186
rect 123 98 126 132
rect 160 98 164 132
rect 123 82 164 98
rect 198 136 280 152
rect 198 102 222 136
rect 256 102 280 136
rect 198 17 280 102
rect 314 136 380 186
rect 314 102 330 136
rect 364 102 380 136
rect 314 86 380 102
rect 414 230 480 236
rect 414 196 430 230
rect 464 196 480 230
rect 414 152 480 196
rect 414 118 430 152
rect 464 118 480 152
rect 414 17 480 118
rect 514 85 548 290
rect 777 256 811 390
rect 1036 358 1070 390
rect 888 344 1070 358
rect 888 310 1020 344
rect 1054 310 1070 344
rect 888 294 1070 310
rect 1127 340 1223 356
rect 1127 306 1143 340
rect 1177 306 1223 340
rect 1127 290 1223 306
rect 1285 354 1319 390
rect 1285 338 1365 354
rect 1285 304 1315 338
rect 1349 304 1365 338
rect 1285 288 1365 304
rect 1413 340 1607 356
rect 1413 306 1429 340
rect 1463 306 1513 340
rect 1547 306 1607 340
rect 1413 290 1607 306
rect 684 253 1226 256
rect 582 226 648 242
rect 582 192 598 226
rect 632 192 648 226
rect 684 219 700 253
rect 734 237 1226 253
rect 734 222 1176 237
rect 734 219 750 222
rect 582 185 648 192
rect 1160 203 1176 222
rect 1210 203 1226 237
rect 870 186 951 188
rect 582 158 786 185
rect 582 124 598 158
rect 632 151 786 158
rect 820 151 836 185
rect 870 152 886 186
rect 920 152 951 186
rect 870 151 951 152
rect 632 124 648 151
rect 582 119 648 124
rect 817 101 883 117
rect 817 85 833 101
rect 514 67 833 85
rect 867 67 883 101
rect 514 51 883 67
rect 917 17 951 151
rect 988 170 1038 188
rect 988 136 1004 170
rect 988 85 1038 136
rect 1074 170 1124 188
rect 1160 187 1226 203
rect 1262 238 1312 254
rect 1296 204 1312 238
rect 1074 136 1090 170
rect 1262 169 1312 204
rect 1124 136 1262 153
rect 1074 135 1262 136
rect 1296 135 1312 169
rect 1074 119 1312 135
rect 1348 238 1609 254
rect 1348 204 1364 238
rect 1398 220 1559 238
rect 1348 168 1398 204
rect 1543 204 1559 220
rect 1593 204 1609 238
rect 1348 134 1364 168
rect 1348 85 1398 134
rect 988 51 1398 85
rect 1438 168 1509 184
rect 1438 134 1456 168
rect 1490 134 1509 168
rect 1438 17 1509 134
rect 1543 168 1609 204
rect 1543 134 1559 168
rect 1593 134 1609 168
rect 1543 118 1609 134
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a32o_4
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 5 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1632 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3712628
string GDS_START 3699320
<< end >>
