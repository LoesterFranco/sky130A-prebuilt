magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1958 704
<< pwell >>
rect 0 0 1920 49
<< scpmos >>
rect 116 387 146 587
rect 235 387 265 587
rect 342 419 372 587
rect 443 419 473 547
rect 533 419 563 547
rect 640 379 670 547
rect 963 368 993 592
rect 1165 424 1195 592
rect 1317 424 1347 592
rect 1535 368 1565 496
rect 1714 368 1744 592
rect 1804 368 1834 592
<< nmoslvt >>
rect 84 134 114 262
rect 250 134 280 262
rect 386 113 416 241
rect 486 157 516 241
rect 620 113 650 241
rect 738 125 768 253
rect 972 74 1002 222
rect 1216 107 1246 235
rect 1352 121 1382 249
rect 1600 78 1630 162
rect 1716 78 1746 226
rect 1802 78 1832 226
<< ndiff >>
rect 27 248 84 262
rect 27 214 39 248
rect 73 214 84 248
rect 27 180 84 214
rect 27 146 39 180
rect 73 146 84 180
rect 27 134 84 146
rect 114 134 250 262
rect 280 250 337 262
rect 280 216 291 250
rect 325 241 337 250
rect 665 241 738 253
rect 325 216 386 241
rect 280 134 386 216
rect 129 82 235 134
rect 336 113 386 134
rect 416 229 486 241
rect 416 195 427 229
rect 461 195 486 229
rect 416 159 486 195
rect 416 125 427 159
rect 461 157 486 159
rect 516 216 620 241
rect 516 182 541 216
rect 575 182 620 216
rect 516 157 620 182
rect 461 125 471 157
rect 416 113 471 125
rect 531 113 620 157
rect 650 207 677 241
rect 711 207 738 241
rect 650 159 738 207
rect 650 125 677 159
rect 711 125 738 159
rect 768 237 857 253
rect 768 203 813 237
rect 847 203 857 237
rect 768 125 857 203
rect 650 113 723 125
rect 129 48 165 82
rect 199 48 235 82
rect 129 36 235 48
rect 1295 237 1352 249
rect 1295 235 1307 237
rect 917 177 972 222
rect 917 143 927 177
rect 961 143 972 177
rect 917 74 972 143
rect 1002 85 1107 222
rect 1161 153 1216 235
rect 1161 119 1171 153
rect 1205 119 1216 153
rect 1161 107 1216 119
rect 1246 203 1307 235
rect 1341 203 1352 237
rect 1246 121 1352 203
rect 1382 169 1449 249
rect 1645 214 1716 226
rect 1382 135 1398 169
rect 1432 135 1449 169
rect 1645 180 1657 214
rect 1691 180 1716 214
rect 1645 162 1716 180
rect 1382 121 1449 135
rect 1543 137 1600 162
rect 1246 107 1296 121
rect 1002 74 1063 85
rect 1017 51 1063 74
rect 1097 51 1107 85
rect 1543 103 1555 137
rect 1589 103 1600 137
rect 1543 78 1600 103
rect 1630 124 1716 162
rect 1630 90 1657 124
rect 1691 90 1716 124
rect 1630 78 1716 90
rect 1746 214 1802 226
rect 1746 180 1757 214
rect 1791 180 1802 214
rect 1746 124 1802 180
rect 1746 90 1757 124
rect 1791 90 1802 124
rect 1746 78 1802 90
rect 1832 214 1889 226
rect 1832 180 1843 214
rect 1877 180 1889 214
rect 1832 124 1889 180
rect 1832 90 1843 124
rect 1877 90 1889 124
rect 1832 78 1889 90
rect 1017 39 1107 51
<< pdiff >>
rect 57 575 116 587
rect 57 541 69 575
rect 103 541 116 575
rect 57 502 116 541
rect 57 468 69 502
rect 103 468 116 502
rect 57 387 116 468
rect 146 575 235 587
rect 146 541 169 575
rect 203 541 235 575
rect 146 502 235 541
rect 146 468 169 502
rect 203 468 235 502
rect 146 387 235 468
rect 265 575 342 587
rect 265 541 278 575
rect 312 541 342 575
rect 265 465 342 541
rect 265 431 278 465
rect 312 431 342 465
rect 265 419 342 431
rect 372 547 425 587
rect 372 533 443 547
rect 372 499 386 533
rect 420 499 443 533
rect 372 465 443 499
rect 372 431 386 465
rect 420 431 443 465
rect 372 419 443 431
rect 473 472 533 547
rect 473 438 486 472
rect 520 438 533 472
rect 473 419 533 438
rect 563 444 640 547
rect 563 419 593 444
rect 265 387 324 419
rect 581 410 593 419
rect 627 410 640 444
rect 581 379 640 410
rect 670 535 802 547
rect 670 501 745 535
rect 779 501 802 535
rect 670 431 802 501
rect 670 397 745 431
rect 779 397 802 431
rect 670 379 802 397
rect 904 580 963 592
rect 904 546 916 580
rect 950 546 963 580
rect 904 497 963 546
rect 904 463 916 497
rect 950 463 963 497
rect 904 414 963 463
rect 904 380 916 414
rect 950 380 963 414
rect 904 368 963 380
rect 993 580 1052 592
rect 993 546 1006 580
rect 1040 546 1052 580
rect 993 497 1052 546
rect 993 463 1006 497
rect 1040 463 1052 497
rect 993 414 1052 463
rect 1106 580 1165 592
rect 1106 546 1118 580
rect 1152 546 1165 580
rect 1106 470 1165 546
rect 1106 436 1118 470
rect 1152 436 1165 470
rect 1106 424 1165 436
rect 1195 504 1317 592
rect 1195 470 1270 504
rect 1304 470 1317 504
rect 1195 424 1317 470
rect 1347 504 1406 592
rect 1583 582 1714 592
rect 1583 580 1667 582
rect 1583 546 1595 580
rect 1629 548 1667 580
rect 1701 548 1714 582
rect 1629 546 1714 548
rect 1347 470 1360 504
rect 1394 470 1406 504
rect 1583 514 1714 546
rect 1583 497 1667 514
rect 1583 496 1595 497
rect 1347 424 1406 470
rect 1460 478 1535 496
rect 1460 444 1472 478
rect 1506 444 1535 478
rect 993 380 1006 414
rect 1040 380 1052 414
rect 993 368 1052 380
rect 1460 368 1535 444
rect 1565 463 1595 496
rect 1629 480 1667 497
rect 1701 480 1714 514
rect 1629 463 1714 480
rect 1565 414 1714 463
rect 1565 380 1595 414
rect 1629 380 1714 414
rect 1565 368 1714 380
rect 1744 580 1804 592
rect 1744 546 1757 580
rect 1791 546 1804 580
rect 1744 497 1804 546
rect 1744 463 1757 497
rect 1791 463 1804 497
rect 1744 414 1804 463
rect 1744 380 1757 414
rect 1791 380 1804 414
rect 1744 368 1804 380
rect 1834 580 1893 592
rect 1834 546 1847 580
rect 1881 546 1893 580
rect 1834 497 1893 546
rect 1834 463 1847 497
rect 1881 463 1893 497
rect 1834 414 1893 463
rect 1834 380 1847 414
rect 1881 380 1893 414
rect 1834 368 1893 380
<< ndiffc >>
rect 39 214 73 248
rect 39 146 73 180
rect 291 216 325 250
rect 427 195 461 229
rect 427 125 461 159
rect 541 182 575 216
rect 677 207 711 241
rect 677 125 711 159
rect 813 203 847 237
rect 165 48 199 82
rect 927 143 961 177
rect 1171 119 1205 153
rect 1307 203 1341 237
rect 1398 135 1432 169
rect 1657 180 1691 214
rect 1063 51 1097 85
rect 1555 103 1589 137
rect 1657 90 1691 124
rect 1757 180 1791 214
rect 1757 90 1791 124
rect 1843 180 1877 214
rect 1843 90 1877 124
<< pdiffc >>
rect 69 541 103 575
rect 69 468 103 502
rect 169 541 203 575
rect 169 468 203 502
rect 278 541 312 575
rect 278 431 312 465
rect 386 499 420 533
rect 386 431 420 465
rect 486 438 520 472
rect 593 410 627 444
rect 745 501 779 535
rect 745 397 779 431
rect 916 546 950 580
rect 916 463 950 497
rect 916 380 950 414
rect 1006 546 1040 580
rect 1006 463 1040 497
rect 1118 546 1152 580
rect 1118 436 1152 470
rect 1270 470 1304 504
rect 1595 546 1629 580
rect 1667 548 1701 582
rect 1360 470 1394 504
rect 1472 444 1506 478
rect 1006 380 1040 414
rect 1595 463 1629 497
rect 1667 480 1701 514
rect 1595 380 1629 414
rect 1757 546 1791 580
rect 1757 463 1791 497
rect 1757 380 1791 414
rect 1847 546 1881 580
rect 1847 463 1881 497
rect 1847 380 1881 414
<< poly >>
rect 339 615 889 645
rect 116 587 146 613
rect 235 587 265 613
rect 339 602 375 615
rect 342 587 372 602
rect 443 547 473 573
rect 530 562 566 615
rect 533 547 563 562
rect 640 547 670 573
rect 342 393 372 419
rect 443 404 473 419
rect 116 372 146 387
rect 235 372 265 387
rect 113 355 149 372
rect 83 339 149 355
rect 232 350 268 372
rect 83 305 99 339
rect 133 305 149 339
rect 83 289 149 305
rect 191 334 280 350
rect 191 300 207 334
rect 241 300 280 334
rect 440 345 476 404
rect 533 393 563 419
rect 640 364 670 379
rect 637 345 673 364
rect 738 345 811 347
rect 440 331 811 345
rect 440 315 761 331
rect 84 262 114 289
rect 191 284 280 300
rect 250 262 280 284
rect 386 241 416 267
rect 486 241 516 315
rect 738 297 761 315
rect 795 297 811 331
rect 738 281 811 297
rect 859 304 889 615
rect 963 592 993 618
rect 1165 592 1195 618
rect 1317 592 1347 618
rect 1714 592 1744 618
rect 1804 592 1834 618
rect 1535 496 1565 522
rect 1165 409 1195 424
rect 1317 409 1347 424
rect 1162 379 1246 409
rect 963 353 993 368
rect 960 310 996 353
rect 1216 337 1246 379
rect 1170 321 1246 337
rect 620 241 650 267
rect 738 253 768 281
rect 859 274 902 304
rect 960 294 1050 310
rect 960 274 1000 294
rect 872 260 1000 274
rect 1034 260 1050 294
rect 1170 287 1186 321
rect 1220 287 1246 321
rect 1314 337 1350 409
rect 1535 353 1565 368
rect 1714 353 1744 368
rect 1804 353 1834 368
rect 1314 321 1428 337
rect 1314 307 1378 321
rect 1170 271 1246 287
rect 84 108 114 134
rect 250 108 280 134
rect 486 131 516 157
rect 872 244 1050 260
rect 386 51 416 113
rect 620 51 650 113
rect 738 99 768 125
rect 872 51 902 244
rect 972 222 1002 244
rect 1216 235 1246 271
rect 1352 287 1378 307
rect 1412 301 1428 321
rect 1532 301 1568 353
rect 1711 330 1747 353
rect 1639 314 1747 330
rect 1412 287 1562 301
rect 1352 271 1562 287
rect 1352 249 1382 271
rect 1532 207 1562 271
rect 1639 280 1655 314
rect 1689 294 1747 314
rect 1801 294 1837 353
rect 1689 280 1837 294
rect 1639 264 1837 280
rect 1716 226 1746 264
rect 1802 226 1832 264
rect 1532 177 1630 207
rect 1600 162 1630 177
rect 386 21 902 51
rect 972 48 1002 74
rect 1216 81 1246 107
rect 1352 95 1382 121
rect 1600 52 1630 78
rect 1716 52 1746 78
rect 1802 52 1832 78
<< polycont >>
rect 99 305 133 339
rect 207 300 241 334
rect 761 297 795 331
rect 1000 260 1034 294
rect 1186 287 1220 321
rect 1378 287 1412 321
rect 1655 280 1689 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 17 575 119 591
rect 17 541 69 575
rect 103 541 119 575
rect 17 502 119 541
rect 17 468 69 502
rect 103 468 119 502
rect 17 452 119 468
rect 153 575 219 649
rect 153 541 169 575
rect 203 541 219 575
rect 153 502 219 541
rect 153 468 169 502
rect 203 468 219 502
rect 153 452 219 468
rect 262 581 779 615
rect 262 575 328 581
rect 262 541 278 575
rect 312 541 328 575
rect 745 551 779 581
rect 916 580 950 596
rect 262 465 328 541
rect 17 255 51 452
rect 262 431 278 465
rect 312 431 328 465
rect 262 418 328 431
rect 85 415 328 418
rect 370 533 711 547
rect 370 499 386 533
rect 420 513 711 533
rect 420 499 436 513
rect 370 465 436 499
rect 370 431 386 465
rect 420 431 436 465
rect 370 415 436 431
rect 470 472 536 479
rect 470 438 486 472
rect 520 438 536 472
rect 85 384 325 415
rect 85 339 149 384
rect 85 305 99 339
rect 133 305 149 339
rect 85 289 149 305
rect 191 334 257 350
rect 191 300 207 334
rect 241 300 257 334
rect 17 248 89 255
rect 17 214 39 248
rect 73 214 89 248
rect 191 236 257 300
rect 291 250 325 384
rect 470 313 536 438
rect 577 444 643 479
rect 577 410 593 444
rect 627 424 643 444
rect 577 390 607 410
rect 641 390 643 424
rect 577 375 643 390
rect 17 180 89 214
rect 291 200 325 216
rect 359 279 536 313
rect 17 146 39 180
rect 73 166 89 180
rect 359 166 393 279
rect 502 245 536 279
rect 73 146 393 166
rect 17 132 393 146
rect 427 229 461 245
rect 427 159 461 195
rect 17 130 89 132
rect 502 216 575 245
rect 502 182 541 216
rect 502 153 575 182
rect 427 119 461 125
rect 609 119 643 375
rect 125 82 239 98
rect 427 85 643 119
rect 677 241 711 513
rect 745 535 879 551
rect 779 501 879 535
rect 745 431 879 501
rect 779 397 879 431
rect 745 381 879 397
rect 677 159 711 207
rect 677 85 711 125
rect 745 331 811 347
rect 745 297 761 331
rect 795 297 811 331
rect 745 287 811 297
rect 745 153 779 287
rect 845 253 879 381
rect 813 237 879 253
rect 847 203 879 237
rect 813 187 879 203
rect 916 497 950 546
rect 916 414 950 463
rect 916 202 950 380
rect 990 580 1040 649
rect 990 546 1006 580
rect 990 497 1040 546
rect 990 463 1006 497
rect 990 414 1040 463
rect 990 380 1006 414
rect 1081 580 1168 596
rect 1081 546 1118 580
rect 1152 546 1168 580
rect 1081 470 1168 546
rect 1081 436 1118 470
rect 1152 436 1168 470
rect 1081 424 1168 436
rect 1081 390 1087 424
rect 1121 390 1168 424
rect 1081 384 1168 390
rect 1202 581 1490 615
rect 990 364 1040 380
rect 984 294 1050 310
rect 984 260 1000 294
rect 1034 260 1050 294
rect 984 236 1050 260
rect 1102 237 1136 384
rect 1202 337 1236 581
rect 1170 321 1236 337
rect 1170 287 1186 321
rect 1220 287 1236 321
rect 1170 271 1236 287
rect 1270 504 1320 540
rect 1304 470 1320 504
rect 1270 424 1320 470
rect 1270 390 1279 424
rect 1313 390 1320 424
rect 1270 305 1320 390
rect 1357 504 1410 538
rect 1357 470 1360 504
rect 1394 470 1410 504
rect 1357 405 1410 470
rect 1456 500 1490 581
rect 1595 582 1706 649
rect 1595 580 1667 582
rect 1629 548 1667 580
rect 1701 548 1706 582
rect 1629 546 1706 548
rect 1595 514 1706 546
rect 1456 478 1561 500
rect 1456 444 1472 478
rect 1506 444 1561 478
rect 1456 439 1561 444
rect 1357 371 1493 405
rect 1375 321 1425 337
rect 1270 271 1341 305
rect 1307 237 1341 271
rect 1102 203 1273 237
rect 916 177 961 202
rect 916 153 927 177
rect 745 143 927 153
rect 745 119 961 143
rect 995 153 1205 169
rect 995 135 1171 153
rect 995 85 1029 135
rect 1155 119 1171 135
rect 1239 153 1273 203
rect 1375 287 1378 321
rect 1412 287 1425 321
rect 1375 236 1425 287
rect 1459 253 1493 371
rect 1527 321 1561 439
rect 1595 497 1667 514
rect 1629 480 1667 497
rect 1701 480 1706 514
rect 1629 464 1706 480
rect 1741 580 1807 596
rect 1741 546 1757 580
rect 1791 546 1807 580
rect 1741 497 1807 546
rect 1595 414 1629 463
rect 1741 463 1757 497
rect 1791 463 1807 497
rect 1595 364 1629 380
rect 1663 424 1705 430
rect 1697 390 1705 424
rect 1663 330 1705 390
rect 1527 287 1605 321
rect 1459 219 1521 253
rect 1307 187 1341 203
rect 1377 169 1453 185
rect 1377 153 1398 169
rect 1239 135 1398 153
rect 1432 135 1453 169
rect 1239 119 1453 135
rect 125 48 165 82
rect 199 48 239 82
rect 677 51 1029 85
rect 1063 85 1113 101
rect 1097 51 1113 85
rect 1155 85 1205 119
rect 1487 85 1521 219
rect 1155 51 1521 85
rect 1555 137 1605 287
rect 1639 314 1705 330
rect 1639 280 1655 314
rect 1689 280 1705 314
rect 1639 264 1705 280
rect 1741 414 1807 463
rect 1741 380 1757 414
rect 1791 380 1807 414
rect 1589 103 1605 137
rect 1555 74 1605 103
rect 1641 214 1707 230
rect 1641 180 1657 214
rect 1691 180 1707 214
rect 1641 124 1707 180
rect 1641 90 1657 124
rect 1691 90 1707 124
rect 125 17 239 48
rect 1063 17 1113 51
rect 1641 17 1707 90
rect 1741 214 1807 380
rect 1847 580 1897 649
rect 1881 546 1897 580
rect 1847 497 1897 546
rect 1881 463 1897 497
rect 1847 414 1897 463
rect 1881 380 1897 414
rect 1847 364 1897 380
rect 1741 180 1757 214
rect 1791 180 1807 214
rect 1741 124 1807 180
rect 1741 90 1757 124
rect 1791 90 1807 124
rect 1741 74 1807 90
rect 1843 214 1893 230
rect 1877 180 1893 214
rect 1843 124 1893 180
rect 1877 90 1893 124
rect 1843 17 1893 90
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 607 410 627 424
rect 627 410 641 424
rect 607 390 641 410
rect 1087 390 1121 424
rect 1279 390 1313 424
rect 1663 390 1697 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 595 424 653 430
rect 595 390 607 424
rect 641 421 653 424
rect 1075 424 1133 430
rect 1075 421 1087 424
rect 641 393 1087 421
rect 641 390 653 393
rect 595 384 653 390
rect 1075 390 1087 393
rect 1121 390 1133 424
rect 1075 384 1133 390
rect 1267 424 1325 430
rect 1267 390 1279 424
rect 1313 421 1325 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 1313 393 1663 421
rect 1313 390 1325 393
rect 1267 384 1325 390
rect 1651 390 1663 393
rect 1697 390 1709 424
rect 1651 384 1709 390
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xor3_2
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 991 242 1025 276 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 1759 94 1793 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 168 1793 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 242 1793 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 316 1793 350 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 390 1793 424 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 464 1793 498 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1759 538 1793 572 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1920 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 600172
string GDS_START 585588
<< end >>
