magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 0 0 1056 49
<< scnmos >>
rect 81 74 111 158
rect 252 74 288 158
rect 513 74 549 158
rect 799 74 835 158
rect 927 74 957 158
<< pmoshvt >>
rect 84 368 114 592
rect 239 392 289 592
rect 499 392 549 592
rect 784 392 834 592
rect 929 368 959 592
<< ndiff >>
rect 28 133 81 158
rect 28 99 36 133
rect 70 99 81 133
rect 28 74 81 99
rect 111 130 252 158
rect 111 96 133 130
rect 167 96 252 130
rect 111 74 252 96
rect 288 133 341 158
rect 288 99 299 133
rect 333 99 341 133
rect 288 74 341 99
rect 395 133 513 158
rect 395 99 404 133
rect 438 99 513 133
rect 395 74 513 99
rect 549 133 602 158
rect 549 99 560 133
rect 594 99 602 133
rect 549 74 602 99
rect 682 130 799 158
rect 682 96 690 130
rect 724 96 799 130
rect 682 74 799 96
rect 835 134 927 158
rect 835 100 882 134
rect 916 100 927 134
rect 835 74 927 100
rect 957 135 1010 158
rect 957 101 968 135
rect 1002 101 1010 135
rect 957 74 1010 101
<< pdiff >>
rect 28 529 84 592
rect 28 495 36 529
rect 70 495 84 529
rect 28 440 84 495
rect 28 406 36 440
rect 70 406 84 440
rect 28 368 84 406
rect 114 584 239 592
rect 114 550 131 584
rect 165 550 239 584
rect 114 510 239 550
rect 114 476 131 510
rect 165 476 239 510
rect 114 392 239 476
rect 289 580 341 592
rect 289 546 299 580
rect 333 546 341 580
rect 289 509 341 546
rect 289 475 299 509
rect 333 475 341 509
rect 289 438 341 475
rect 289 404 299 438
rect 333 404 341 438
rect 289 392 341 404
rect 395 580 499 592
rect 395 546 403 580
rect 437 546 499 580
rect 395 509 499 546
rect 395 475 403 509
rect 437 475 499 509
rect 395 438 499 475
rect 395 404 403 438
rect 437 404 499 438
rect 395 392 499 404
rect 549 580 602 592
rect 549 546 560 580
rect 594 546 602 580
rect 549 509 602 546
rect 549 475 560 509
rect 594 475 602 509
rect 549 438 602 475
rect 549 404 560 438
rect 594 404 602 438
rect 549 392 602 404
rect 682 580 784 592
rect 682 546 690 580
rect 724 546 784 580
rect 682 509 784 546
rect 682 475 690 509
rect 724 475 784 509
rect 682 438 784 475
rect 682 404 690 438
rect 724 404 784 438
rect 682 392 784 404
rect 834 579 929 592
rect 834 545 882 579
rect 916 545 929 579
rect 834 500 929 545
rect 834 466 882 500
rect 916 466 929 500
rect 834 414 929 466
rect 834 392 882 414
rect 114 368 167 392
rect 874 380 882 392
rect 916 380 929 414
rect 874 368 929 380
rect 959 579 1015 592
rect 959 545 973 579
rect 1007 545 1015 579
rect 959 507 1015 545
rect 959 473 973 507
rect 1007 473 1015 507
rect 959 430 1015 473
rect 959 396 973 430
rect 1007 396 1015 430
rect 959 368 1015 396
<< ndiffc >>
rect 36 99 70 133
rect 133 96 167 130
rect 299 99 333 133
rect 404 99 438 133
rect 560 99 594 133
rect 690 96 724 130
rect 882 100 916 134
rect 968 101 1002 135
<< pdiffc >>
rect 36 495 70 529
rect 36 406 70 440
rect 131 550 165 584
rect 131 476 165 510
rect 299 546 333 580
rect 299 475 333 509
rect 299 404 333 438
rect 403 546 437 580
rect 403 475 437 509
rect 403 404 437 438
rect 560 546 594 580
rect 560 475 594 509
rect 560 404 594 438
rect 690 546 724 580
rect 690 475 724 509
rect 690 404 724 438
rect 882 545 916 579
rect 882 466 916 500
rect 882 380 916 414
rect 973 545 1007 579
rect 973 473 1007 507
rect 973 396 1007 430
<< poly >>
rect 84 592 114 618
rect 239 592 289 618
rect 499 592 549 618
rect 784 592 834 618
rect 929 592 959 618
rect 84 353 114 368
rect 81 304 117 353
rect 81 288 147 304
rect 239 292 289 392
rect 499 294 549 392
rect 784 294 834 392
rect 929 353 959 368
rect 926 325 962 353
rect 81 254 97 288
rect 131 254 147 288
rect 81 238 147 254
rect 189 276 289 292
rect 189 242 211 276
rect 245 242 289 276
rect 81 158 111 238
rect 189 226 289 242
rect 449 278 549 294
rect 449 244 468 278
rect 502 244 549 278
rect 449 228 549 244
rect 734 278 834 294
rect 734 244 751 278
rect 785 259 834 278
rect 901 309 967 325
rect 901 275 917 309
rect 951 275 967 309
rect 901 259 967 275
rect 785 244 835 259
rect 734 228 835 244
rect 252 158 288 226
rect 513 158 549 228
rect 799 158 835 228
rect 927 158 957 259
rect 81 48 111 74
rect 252 48 288 74
rect 513 48 549 74
rect 799 48 835 74
rect 927 48 957 74
<< polycont >>
rect 97 254 131 288
rect 211 242 245 276
rect 468 244 502 278
rect 751 244 785 278
rect 917 275 951 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 115 584 181 649
rect 115 550 131 584
rect 165 550 181 584
rect 383 580 453 649
rect 19 529 80 545
rect 19 495 36 529
rect 70 495 80 529
rect 19 441 80 495
rect 115 510 181 550
rect 283 546 299 580
rect 333 546 349 580
rect 283 530 349 546
rect 115 476 131 510
rect 165 476 181 510
rect 295 509 349 530
rect 295 475 299 509
rect 333 475 349 509
rect 19 440 261 441
rect 19 406 36 440
rect 70 406 261 440
rect 20 288 146 372
rect 20 254 97 288
rect 131 254 146 288
rect 20 238 146 254
rect 195 276 261 406
rect 195 242 211 276
rect 245 242 261 276
rect 195 204 261 242
rect 19 164 261 204
rect 295 438 349 475
rect 295 404 299 438
rect 333 404 349 438
rect 295 294 349 404
rect 383 546 403 580
rect 437 546 453 580
rect 383 509 453 546
rect 383 475 403 509
rect 437 475 453 509
rect 383 438 453 475
rect 383 404 403 438
rect 437 404 453 438
rect 383 388 453 404
rect 560 580 594 596
rect 560 509 594 546
rect 560 438 594 475
rect 295 278 502 294
rect 295 244 468 278
rect 295 228 502 244
rect 560 278 594 404
rect 683 580 731 596
rect 683 546 690 580
rect 724 546 731 580
rect 683 509 731 546
rect 683 475 690 509
rect 724 475 731 509
rect 683 438 731 475
rect 683 404 690 438
rect 724 404 731 438
rect 683 346 731 404
rect 866 579 932 649
rect 866 545 882 579
rect 916 545 932 579
rect 866 500 932 545
rect 866 466 882 500
rect 916 466 932 500
rect 866 414 932 466
rect 866 380 882 414
rect 916 380 932 414
rect 966 579 1038 612
rect 966 545 973 579
rect 1007 545 1038 579
rect 966 507 1038 545
rect 966 473 973 507
rect 1007 473 1038 507
rect 966 430 1038 473
rect 966 396 973 430
rect 1007 396 1038 430
rect 966 380 1038 396
rect 683 312 951 346
rect 906 309 951 312
rect 560 244 751 278
rect 785 244 801 278
rect 906 275 917 309
rect 19 133 82 164
rect 19 99 36 133
rect 70 99 82 133
rect 295 133 344 228
rect 19 61 82 99
rect 117 96 133 130
rect 167 96 183 130
rect 117 17 183 96
rect 295 99 299 133
rect 333 99 344 133
rect 295 61 344 99
rect 383 133 453 149
rect 383 99 404 133
rect 438 99 453 133
rect 383 17 453 99
rect 560 133 594 244
rect 906 210 951 275
rect 560 83 594 99
rect 674 185 951 210
rect 674 176 940 185
rect 674 130 740 176
rect 985 151 1038 380
rect 966 135 1038 151
rect 674 96 690 130
rect 724 96 740 130
rect 674 80 740 96
rect 866 100 882 134
rect 916 100 932 134
rect 866 17 932 100
rect 966 101 968 135
rect 1002 101 1038 135
rect 966 71 1038 101
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 clkdlyinv5sd2_1
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 990 464 1024 498 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 990 390 1024 424 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 990 168 1024 202 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 990 94 1024 128 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 990 242 1024 276 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel corelocali s 990 538 1024 572 0 FreeSans 200 0 0 0 Y
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 1056 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3370736
string GDS_START 3362764
<< end >>
