magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scnmos >>
rect 85 138 115 248
rect 188 100 218 248
rect 274 100 304 248
rect 421 120 451 248
rect 548 136 578 264
rect 656 136 686 264
rect 744 136 774 264
rect 846 91 876 201
<< pmoshvt >>
rect 84 424 114 592
rect 185 368 215 592
rect 275 368 305 592
rect 473 392 503 592
rect 557 392 587 592
rect 659 392 689 592
rect 737 392 767 592
rect 845 392 875 560
<< ndiff >>
rect 466 248 548 264
rect 28 202 85 248
rect 28 168 40 202
rect 74 168 85 202
rect 28 138 85 168
rect 115 149 188 248
rect 115 138 142 149
rect 130 115 142 138
rect 176 115 188 149
rect 130 100 188 115
rect 218 220 274 248
rect 218 186 229 220
rect 263 186 274 220
rect 218 146 274 186
rect 218 112 229 146
rect 263 112 274 146
rect 218 100 274 112
rect 304 175 421 248
rect 304 141 347 175
rect 381 141 421 175
rect 304 120 421 141
rect 451 236 548 248
rect 451 202 478 236
rect 512 202 548 236
rect 451 166 548 202
rect 451 132 478 166
rect 512 136 548 166
rect 578 187 656 264
rect 578 153 589 187
rect 623 153 656 187
rect 578 136 656 153
rect 686 231 744 264
rect 686 197 697 231
rect 731 197 744 231
rect 686 136 744 197
rect 774 201 824 264
rect 774 139 846 201
rect 774 136 801 139
rect 512 132 524 136
rect 451 120 524 132
rect 304 100 354 120
rect 789 105 801 136
rect 835 105 846 139
rect 789 91 846 105
rect 876 163 933 201
rect 876 129 887 163
rect 921 129 933 163
rect 876 91 933 129
<< pdiff >>
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 470 84 546
rect 27 436 37 470
rect 71 436 84 470
rect 27 424 84 436
rect 114 576 185 592
rect 114 542 137 576
rect 171 542 185 576
rect 114 424 185 542
rect 132 368 185 424
rect 215 420 275 592
rect 215 386 228 420
rect 262 386 275 420
rect 215 368 275 386
rect 305 576 362 592
rect 305 542 318 576
rect 352 542 362 576
rect 305 368 362 542
rect 416 576 473 592
rect 416 542 426 576
rect 460 542 473 576
rect 416 392 473 542
rect 503 392 557 592
rect 587 392 659 592
rect 689 392 737 592
rect 767 576 826 592
rect 767 542 780 576
rect 814 560 826 576
rect 814 542 845 560
rect 767 496 845 542
rect 767 462 780 496
rect 814 462 845 496
rect 767 392 845 462
rect 875 548 933 560
rect 875 514 888 548
rect 922 514 933 548
rect 875 440 933 514
rect 875 406 888 440
rect 922 406 933 440
rect 875 392 933 406
<< ndiffc >>
rect 40 168 74 202
rect 142 115 176 149
rect 229 186 263 220
rect 229 112 263 146
rect 347 141 381 175
rect 478 202 512 236
rect 478 132 512 166
rect 589 153 623 187
rect 697 197 731 231
rect 801 105 835 139
rect 887 129 921 163
<< pdiffc >>
rect 37 546 71 580
rect 37 436 71 470
rect 137 542 171 576
rect 228 386 262 420
rect 318 542 352 576
rect 426 542 460 576
rect 780 542 814 576
rect 780 462 814 496
rect 888 514 922 548
rect 888 406 922 440
<< poly >>
rect 84 592 114 618
rect 185 592 215 618
rect 275 592 305 618
rect 473 592 503 618
rect 557 592 587 618
rect 659 592 689 618
rect 737 592 767 618
rect 84 409 114 424
rect 81 336 117 409
rect 845 560 875 586
rect 473 377 503 392
rect 557 377 587 392
rect 659 377 689 392
rect 737 377 767 392
rect 845 377 875 392
rect 185 353 215 368
rect 275 353 305 368
rect 470 360 506 377
rect 554 360 590 377
rect 44 320 115 336
rect 44 286 60 320
rect 94 286 115 320
rect 44 270 115 286
rect 182 317 218 353
rect 272 336 308 353
rect 394 344 506 360
rect 272 320 346 336
rect 272 317 296 320
rect 182 286 296 317
rect 330 286 346 320
rect 394 310 410 344
rect 444 310 506 344
rect 394 294 506 310
rect 548 344 614 360
rect 548 310 564 344
rect 598 310 614 344
rect 548 294 614 310
rect 182 270 346 286
rect 85 248 115 270
rect 188 248 218 270
rect 274 248 304 270
rect 421 248 451 294
rect 548 264 578 294
rect 656 279 692 377
rect 734 360 770 377
rect 734 344 800 360
rect 734 310 750 344
rect 784 310 800 344
rect 734 294 800 310
rect 842 326 878 377
rect 842 310 939 326
rect 656 264 686 279
rect 744 264 774 294
rect 842 276 889 310
rect 923 276 939 310
rect 85 112 115 138
rect 842 260 939 276
rect 846 201 876 260
rect 188 74 218 100
rect 274 74 304 100
rect 421 94 451 120
rect 548 110 578 136
rect 656 114 686 136
rect 630 98 696 114
rect 744 110 774 136
rect 630 64 646 98
rect 680 64 696 98
rect 846 65 876 91
rect 630 48 696 64
<< polycont >>
rect 60 286 94 320
rect 296 286 330 320
rect 410 310 444 344
rect 564 310 598 344
rect 750 310 784 344
rect 889 276 923 310
rect 646 64 680 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 21 580 87 596
rect 21 546 37 580
rect 71 546 87 580
rect 21 488 87 546
rect 121 576 187 649
rect 121 542 137 576
rect 171 542 187 576
rect 121 522 187 542
rect 302 576 368 649
rect 302 542 318 576
rect 352 542 368 576
rect 302 522 368 542
rect 410 576 476 596
rect 410 542 426 576
rect 460 556 476 576
rect 764 576 830 649
rect 460 542 521 556
rect 410 522 521 542
rect 21 470 453 488
rect 21 436 37 470
rect 71 454 453 470
rect 71 436 178 454
rect 21 420 178 436
rect 25 320 110 356
rect 25 286 60 320
rect 94 286 110 320
rect 25 270 110 286
rect 144 236 178 420
rect 24 202 178 236
rect 212 386 228 420
rect 262 386 278 420
rect 212 370 278 386
rect 212 236 246 370
rect 394 344 453 454
rect 280 320 346 336
rect 280 286 296 320
rect 330 286 346 320
rect 394 310 410 344
rect 444 310 453 344
rect 394 294 453 310
rect 280 270 346 286
rect 312 260 346 270
rect 487 260 521 522
rect 764 542 780 576
rect 814 542 830 576
rect 764 496 830 542
rect 764 462 780 496
rect 814 462 830 496
rect 872 548 938 564
rect 872 514 888 548
rect 922 514 938 548
rect 872 440 938 514
rect 872 428 888 440
rect 555 406 888 428
rect 922 406 938 440
rect 555 394 938 406
rect 555 344 614 394
rect 819 390 938 394
rect 555 310 564 344
rect 598 310 614 344
rect 555 294 614 310
rect 697 344 785 360
rect 697 310 750 344
rect 784 310 785 344
rect 697 294 785 310
rect 312 236 747 260
rect 212 220 263 236
rect 312 226 478 236
rect 24 168 40 202
rect 74 168 90 202
rect 212 186 229 220
rect 24 134 90 168
rect 126 149 176 168
rect 126 115 142 149
rect 126 17 176 115
rect 212 146 263 186
rect 462 202 478 226
rect 512 231 747 236
rect 512 226 697 231
rect 512 202 528 226
rect 212 112 229 146
rect 212 88 263 112
rect 315 175 407 182
rect 315 141 347 175
rect 381 141 407 175
rect 315 17 407 141
rect 462 166 528 202
rect 681 197 697 226
rect 731 197 747 231
rect 462 132 478 166
rect 512 132 528 166
rect 462 116 528 132
rect 562 187 639 192
rect 562 153 589 187
rect 623 153 639 187
rect 681 168 747 197
rect 819 226 853 390
rect 887 310 939 356
rect 887 276 889 310
rect 923 276 939 310
rect 887 260 939 276
rect 819 192 937 226
rect 887 163 937 192
rect 562 148 639 153
rect 562 17 596 148
rect 785 139 851 158
rect 697 114 743 134
rect 630 98 743 114
rect 630 64 646 98
rect 680 64 743 98
rect 630 51 743 64
rect 785 105 801 139
rect 835 105 851 139
rect 785 17 851 105
rect 921 129 937 163
rect 887 87 937 129
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or4bb_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 960 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 1136710
string GDS_START 1128688
<< end >>
