magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 129 424 163 547
rect 293 424 359 547
rect 947 424 1013 547
rect 1127 424 1193 547
rect 129 390 1195 424
rect 25 286 359 356
rect 409 286 839 356
rect 889 286 1127 356
rect 1161 252 1195 390
rect 1273 270 1703 356
rect 1753 270 2183 356
rect 109 218 1195 252
rect 109 119 175 218
rect 311 119 361 218
rect 495 119 561 218
rect 695 119 761 218
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 581 449 615
rect 23 390 89 581
rect 203 458 253 581
rect 399 492 449 581
rect 489 526 523 649
rect 563 492 629 596
rect 669 526 703 649
rect 745 492 811 596
rect 399 458 811 492
rect 857 581 1693 615
rect 857 458 907 581
rect 1053 458 1087 581
rect 1229 390 1293 581
rect 1327 424 1393 547
rect 1427 458 1493 581
rect 1527 424 1593 547
rect 1627 458 1693 581
rect 1739 458 1789 649
rect 1829 424 1895 596
rect 1929 458 1995 649
rect 2029 424 2095 596
rect 1327 390 2095 424
rect 2135 390 2185 649
rect 23 85 73 226
rect 209 85 275 184
rect 395 85 461 184
rect 595 85 661 184
rect 1266 202 2134 236
rect 1266 184 1334 202
rect 795 150 1334 184
rect 795 85 861 150
rect 23 51 861 85
rect 897 17 963 116
rect 999 66 1065 150
rect 1099 17 1165 116
rect 1199 66 1334 150
rect 1368 17 1434 168
rect 1468 70 1534 202
rect 1568 17 1634 168
rect 1668 70 1734 202
rect 1768 17 1834 168
rect 1868 70 1934 202
rect 1968 17 2034 168
rect 2068 70 2134 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel locali s 1753 270 2183 356 6 A1
port 1 nsew signal input
rlabel locali s 1273 270 1703 356 6 A2
port 2 nsew signal input
rlabel locali s 889 286 1127 356 6 A3
port 3 nsew signal input
rlabel locali s 409 286 839 356 6 B1
port 4 nsew signal input
rlabel locali s 25 286 359 356 6 B2
port 5 nsew signal input
rlabel locali s 1161 252 1195 390 6 Y
port 6 nsew signal output
rlabel locali s 1127 424 1193 547 6 Y
port 6 nsew signal output
rlabel locali s 947 424 1013 547 6 Y
port 6 nsew signal output
rlabel locali s 695 119 761 218 6 Y
port 6 nsew signal output
rlabel locali s 495 119 561 218 6 Y
port 6 nsew signal output
rlabel locali s 311 119 361 218 6 Y
port 6 nsew signal output
rlabel locali s 293 424 359 547 6 Y
port 6 nsew signal output
rlabel locali s 129 424 163 547 6 Y
port 6 nsew signal output
rlabel locali s 129 390 1195 424 6 Y
port 6 nsew signal output
rlabel locali s 109 218 1195 252 6 Y
port 6 nsew signal output
rlabel locali s 109 119 175 218 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -49 2208 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 617 2208 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 642226
string GDS_START 624274
<< end >>
