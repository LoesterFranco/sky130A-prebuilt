magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 24 424 90 596
rect 204 424 270 596
rect 24 390 359 424
rect 25 270 263 356
rect 313 236 359 390
rect 123 202 359 236
rect 123 102 261 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 130 458 164 649
rect 310 458 360 649
rect 23 17 89 168
rect 295 17 361 168
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
rlabel locali s 25 270 263 356 6 A
port 1 nsew signal input
rlabel locali s 313 236 359 390 6 Y
port 2 nsew signal output
rlabel locali s 204 424 270 596 6 Y
port 2 nsew signal output
rlabel locali s 123 202 359 236 6 Y
port 2 nsew signal output
rlabel locali s 123 102 261 202 6 Y
port 2 nsew signal output
rlabel locali s 24 424 90 596 6 Y
port 2 nsew signal output
rlabel locali s 24 390 359 424 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 384 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 384 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 384 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3332200
string GDS_START 3328098
<< end >>
