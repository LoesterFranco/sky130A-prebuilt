magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 29 149 82 265
rect 383 425 498 493
rect 625 359 718 493
rect 397 153 524 249
rect 648 289 718 359
rect 648 185 808 289
rect 397 61 474 153
rect 648 143 714 185
rect 633 51 714 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 315 80 527
rect 216 426 349 527
rect 126 249 181 381
rect 220 319 267 392
rect 301 391 349 426
rect 301 353 377 391
rect 432 319 470 378
rect 532 358 575 527
rect 220 285 604 319
rect 126 203 293 249
rect 17 17 71 115
rect 126 61 181 203
rect 329 114 363 285
rect 221 61 363 114
rect 558 199 604 285
rect 752 325 805 527
rect 522 17 588 116
rect 752 17 805 149
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 29 149 82 265 6 A_N
port 1 nsew signal input
rlabel locali s 383 425 498 493 6 B
port 2 nsew signal input
rlabel locali s 397 153 524 249 6 C
port 3 nsew signal input
rlabel locali s 397 61 474 153 6 C
port 3 nsew signal input
rlabel locali s 648 289 718 359 6 X
port 4 nsew signal output
rlabel locali s 648 185 808 289 6 X
port 4 nsew signal output
rlabel locali s 648 143 714 185 6 X
port 4 nsew signal output
rlabel locali s 633 51 714 143 6 X
port 4 nsew signal output
rlabel locali s 625 359 718 493 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1544568
string GDS_START 1537716
<< end >>
