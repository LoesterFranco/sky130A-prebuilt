magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 119 367 257 527
rect 194 289 257 367
rect 291 333 357 493
rect 391 367 425 527
rect 459 333 528 493
rect 562 367 596 527
rect 630 333 696 493
rect 730 367 764 527
rect 798 333 864 493
rect 291 289 864 333
rect 904 299 970 527
rect 22 215 88 255
rect 475 181 528 289
rect 631 215 988 255
rect 119 17 158 109
rect 291 127 528 181
rect 646 17 680 109
rect 814 17 862 109
rect 0 -17 1012 17
<< obsli1 >>
rect 18 333 85 493
rect 18 289 156 333
rect 122 255 156 289
rect 122 215 441 255
rect 122 181 156 215
rect 18 143 156 181
rect 18 51 85 143
rect 207 93 257 181
rect 562 143 970 181
rect 562 93 612 143
rect 207 51 612 93
rect 714 51 780 143
rect 904 51 970 143
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< labels >>
rlabel locali s 22 215 88 255 6 A_N
port 1 nsew signal input
rlabel locali s 631 215 988 255 6 B
port 2 nsew signal input
rlabel locali s 798 333 864 493 6 Y
port 3 nsew signal output
rlabel locali s 630 333 696 493 6 Y
port 3 nsew signal output
rlabel locali s 475 181 528 289 6 Y
port 3 nsew signal output
rlabel locali s 459 333 528 493 6 Y
port 3 nsew signal output
rlabel locali s 291 333 357 493 6 Y
port 3 nsew signal output
rlabel locali s 291 289 864 333 6 Y
port 3 nsew signal output
rlabel locali s 291 127 528 181 6 Y
port 3 nsew signal output
rlabel locali s 814 17 862 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 646 17 680 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 119 17 158 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 904 299 970 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 730 367 764 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 562 367 596 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 391 367 425 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 194 289 257 367 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 119 367 257 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1788802
string GDS_START 1779746
<< end >>
