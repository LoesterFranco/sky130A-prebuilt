magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 87 368 117 592
rect 179 368 209 592
rect 277 368 307 592
rect 381 368 411 592
rect 583 368 613 592
rect 673 368 703 592
rect 763 368 793 592
rect 853 368 883 592
rect 943 368 973 592
rect 1033 368 1063 592
<< nmoslvt >>
rect 84 74 114 222
rect 182 74 212 222
rect 280 74 310 222
rect 368 74 398 222
rect 462 74 492 222
rect 554 74 584 222
rect 640 74 670 222
rect 754 74 784 222
rect 952 74 982 222
rect 1038 74 1068 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 136 182 222
rect 114 102 125 136
rect 159 102 182 136
rect 114 74 182 102
rect 212 210 280 222
rect 212 176 223 210
rect 257 176 280 210
rect 212 120 280 176
rect 212 86 223 120
rect 257 86 280 120
rect 212 74 280 86
rect 310 136 368 222
rect 310 102 323 136
rect 357 102 368 136
rect 310 74 368 102
rect 398 210 462 222
rect 398 176 409 210
rect 443 176 462 210
rect 398 120 462 176
rect 398 86 409 120
rect 443 86 462 120
rect 398 74 462 86
rect 492 136 554 222
rect 492 102 509 136
rect 543 102 554 136
rect 492 74 554 102
rect 584 210 640 222
rect 584 176 595 210
rect 629 176 640 210
rect 584 120 640 176
rect 584 86 595 120
rect 629 86 640 120
rect 584 74 640 86
rect 670 136 754 222
rect 670 102 695 136
rect 729 102 754 136
rect 670 74 754 102
rect 784 189 841 222
rect 784 155 795 189
rect 829 155 841 189
rect 784 74 841 155
rect 895 189 952 222
rect 895 155 907 189
rect 941 155 952 189
rect 895 74 952 155
rect 982 131 1038 222
rect 982 97 993 131
rect 1027 97 1038 131
rect 982 74 1038 97
rect 1068 210 1125 222
rect 1068 176 1079 210
rect 1113 176 1125 210
rect 1068 120 1125 176
rect 1068 86 1079 120
rect 1113 86 1125 120
rect 1068 74 1125 86
<< pdiff >>
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 510 87 546
rect 28 476 40 510
rect 74 476 87 510
rect 28 440 87 476
rect 28 406 40 440
rect 74 406 87 440
rect 28 368 87 406
rect 117 580 179 592
rect 117 546 130 580
rect 164 546 179 580
rect 117 508 179 546
rect 117 474 130 508
rect 164 474 179 508
rect 117 368 179 474
rect 209 580 277 592
rect 209 546 230 580
rect 264 546 277 580
rect 209 510 277 546
rect 209 476 230 510
rect 264 476 277 510
rect 209 440 277 476
rect 209 406 230 440
rect 264 406 277 440
rect 209 368 277 406
rect 307 580 381 592
rect 307 546 334 580
rect 368 546 381 580
rect 307 508 381 546
rect 307 474 334 508
rect 368 474 381 508
rect 307 368 381 474
rect 411 531 470 592
rect 411 497 424 531
rect 458 497 470 531
rect 411 440 470 497
rect 411 406 424 440
rect 458 406 470 440
rect 411 368 470 406
rect 524 531 583 592
rect 524 497 536 531
rect 570 497 583 531
rect 524 440 583 497
rect 524 406 536 440
rect 570 406 583 440
rect 524 368 583 406
rect 613 580 673 592
rect 613 546 626 580
rect 660 546 673 580
rect 613 508 673 546
rect 613 474 626 508
rect 660 474 673 508
rect 613 368 673 474
rect 703 580 763 592
rect 703 546 716 580
rect 750 546 763 580
rect 703 510 763 546
rect 703 476 716 510
rect 750 476 763 510
rect 703 440 763 476
rect 703 406 716 440
rect 750 406 763 440
rect 703 368 763 406
rect 793 580 853 592
rect 793 546 806 580
rect 840 546 853 580
rect 793 508 853 546
rect 793 474 806 508
rect 840 474 853 508
rect 793 368 853 474
rect 883 580 943 592
rect 883 546 896 580
rect 930 546 943 580
rect 883 497 943 546
rect 883 463 896 497
rect 930 463 943 497
rect 883 414 943 463
rect 883 380 896 414
rect 930 380 943 414
rect 883 368 943 380
rect 973 580 1033 592
rect 973 546 986 580
rect 1020 546 1033 580
rect 973 508 1033 546
rect 973 474 986 508
rect 1020 474 1033 508
rect 973 368 1033 474
rect 1063 580 1122 592
rect 1063 546 1076 580
rect 1110 546 1122 580
rect 1063 510 1122 546
rect 1063 476 1076 510
rect 1110 476 1122 510
rect 1063 440 1122 476
rect 1063 406 1076 440
rect 1110 406 1122 440
rect 1063 368 1122 406
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 102 159 136
rect 223 176 257 210
rect 223 86 257 120
rect 323 102 357 136
rect 409 176 443 210
rect 409 86 443 120
rect 509 102 543 136
rect 595 176 629 210
rect 595 86 629 120
rect 695 102 729 136
rect 795 155 829 189
rect 907 155 941 189
rect 993 97 1027 131
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 474 164 508
rect 230 546 264 580
rect 230 476 264 510
rect 230 406 264 440
rect 334 546 368 580
rect 334 474 368 508
rect 424 497 458 531
rect 424 406 458 440
rect 536 497 570 531
rect 536 406 570 440
rect 626 546 660 580
rect 626 474 660 508
rect 716 546 750 580
rect 716 476 750 510
rect 716 406 750 440
rect 806 546 840 580
rect 806 474 840 508
rect 896 546 930 580
rect 896 463 930 497
rect 896 380 930 414
rect 986 546 1020 580
rect 986 474 1020 508
rect 1076 546 1110 580
rect 1076 476 1110 510
rect 1076 406 1110 440
<< poly >>
rect 87 592 117 618
rect 179 592 209 618
rect 277 592 307 618
rect 381 592 411 618
rect 583 592 613 618
rect 673 592 703 618
rect 763 592 793 618
rect 853 592 883 618
rect 943 592 973 618
rect 1033 592 1063 618
rect 87 353 117 368
rect 179 353 209 368
rect 277 353 307 368
rect 381 353 411 368
rect 583 353 613 368
rect 673 353 703 368
rect 763 353 793 368
rect 853 353 883 368
rect 943 353 973 368
rect 1033 353 1063 368
rect 84 336 120 353
rect 176 336 212 353
rect 277 336 310 353
rect 378 336 414 353
rect 580 345 616 353
rect 670 345 706 353
rect 84 320 212 336
rect 84 286 100 320
rect 134 286 212 320
rect 84 270 212 286
rect 84 222 114 270
rect 182 222 212 270
rect 280 320 414 336
rect 280 286 296 320
rect 330 286 364 320
rect 398 286 414 320
rect 280 270 414 286
rect 462 320 706 345
rect 760 336 796 353
rect 850 336 886 353
rect 462 286 521 320
rect 555 315 706 320
rect 754 320 886 336
rect 555 286 584 315
rect 462 270 584 286
rect 280 222 310 270
rect 368 222 398 270
rect 462 222 492 270
rect 554 222 584 270
rect 754 286 770 320
rect 804 306 886 320
rect 940 326 976 353
rect 1030 326 1066 353
rect 940 310 1119 326
rect 804 286 820 306
rect 754 267 820 286
rect 640 237 820 267
rect 940 276 1001 310
rect 1035 276 1069 310
rect 1103 276 1119 310
rect 940 260 1119 276
rect 640 222 670 237
rect 754 222 784 237
rect 952 222 982 260
rect 1038 222 1068 260
rect 84 48 114 74
rect 182 48 212 74
rect 280 48 310 74
rect 368 48 398 74
rect 462 48 492 74
rect 554 48 584 74
rect 640 48 670 74
rect 754 48 784 74
rect 952 48 982 74
rect 1038 48 1068 74
<< polycont >>
rect 100 286 134 320
rect 296 286 330 320
rect 364 286 398 320
rect 521 286 555 320
rect 770 286 804 320
rect 1001 276 1035 310
rect 1069 276 1103 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 24 580 90 596
rect 24 546 40 580
rect 74 546 90 580
rect 24 510 90 546
rect 24 476 40 510
rect 74 476 90 510
rect 24 440 90 476
rect 130 580 180 649
rect 164 546 180 580
rect 130 508 180 546
rect 164 474 180 508
rect 130 458 180 474
rect 214 580 280 596
rect 214 546 230 580
rect 264 546 280 580
rect 214 510 280 546
rect 214 476 230 510
rect 264 476 280 510
rect 24 406 40 440
rect 74 424 90 440
rect 214 440 280 476
rect 318 581 660 615
rect 318 580 384 581
rect 318 546 334 580
rect 368 546 384 580
rect 626 580 660 581
rect 318 508 384 546
rect 318 474 334 508
rect 368 474 384 508
rect 318 458 384 474
rect 424 531 474 547
rect 458 497 474 531
rect 214 424 230 440
rect 74 406 230 424
rect 264 424 280 440
rect 424 440 474 497
rect 264 406 424 424
rect 458 406 474 440
rect 24 390 474 406
rect 520 531 586 547
rect 520 497 536 531
rect 570 497 586 531
rect 520 440 586 497
rect 626 508 660 546
rect 626 458 660 474
rect 700 580 750 596
rect 700 546 716 580
rect 700 510 750 546
rect 700 476 716 510
rect 520 406 536 440
rect 570 424 586 440
rect 700 440 750 476
rect 790 580 856 649
rect 790 546 806 580
rect 840 546 856 580
rect 790 508 856 546
rect 790 474 806 508
rect 840 474 856 508
rect 790 458 856 474
rect 896 580 930 596
rect 896 497 930 546
rect 700 424 716 440
rect 570 406 716 424
rect 896 424 930 463
rect 970 580 1020 649
rect 970 546 986 580
rect 970 508 1020 546
rect 970 474 986 508
rect 970 458 1020 474
rect 1060 580 1126 596
rect 1060 546 1076 580
rect 1110 546 1126 580
rect 1060 510 1126 546
rect 1060 476 1076 510
rect 1110 476 1126 510
rect 1060 440 1126 476
rect 1060 424 1076 440
rect 750 414 1076 424
rect 750 406 896 414
rect 520 390 896 406
rect 880 380 896 390
rect 930 406 1076 414
rect 1110 406 1126 440
rect 930 390 1126 406
rect 930 380 946 390
rect 25 320 167 356
rect 25 286 100 320
rect 134 286 167 320
rect 25 270 167 286
rect 217 320 455 356
rect 217 286 296 320
rect 330 286 364 320
rect 398 286 455 320
rect 217 270 455 286
rect 505 320 647 356
rect 505 286 521 320
rect 555 286 647 320
rect 505 270 647 286
rect 697 320 839 356
rect 697 286 770 320
rect 804 286 839 320
rect 697 270 839 286
rect 23 210 845 236
rect 23 176 39 210
rect 73 202 223 210
rect 23 120 73 176
rect 257 202 409 210
rect 257 176 273 202
rect 23 86 39 120
rect 23 70 73 86
rect 109 136 175 168
rect 109 102 125 136
rect 159 102 175 136
rect 109 17 175 102
rect 223 120 273 176
rect 443 202 595 210
rect 443 176 459 202
rect 257 86 273 120
rect 223 70 273 86
rect 307 136 373 168
rect 307 102 323 136
rect 357 102 373 136
rect 307 17 373 102
rect 409 120 459 176
rect 629 202 845 210
rect 629 176 645 202
rect 443 86 459 120
rect 409 70 459 86
rect 493 136 559 168
rect 493 102 509 136
rect 543 102 559 136
rect 493 17 559 102
rect 595 120 645 176
rect 779 189 845 202
rect 629 86 645 120
rect 595 70 645 86
rect 679 136 745 168
rect 679 102 695 136
rect 729 102 745 136
rect 779 155 795 189
rect 829 155 845 189
rect 779 119 845 155
rect 880 226 946 380
rect 985 310 1127 356
rect 985 276 1001 310
rect 1035 276 1069 310
rect 1103 276 1127 310
rect 985 260 1127 276
rect 880 210 1129 226
rect 880 192 1079 210
rect 880 189 941 192
rect 880 155 907 189
rect 1113 176 1129 210
rect 880 119 941 155
rect 977 131 1043 158
rect 679 85 745 102
rect 977 97 993 131
rect 1027 97 1043 131
rect 977 85 1043 97
rect 679 51 1043 85
rect 1079 120 1129 176
rect 1113 86 1129 120
rect 1079 70 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o311ai_2
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C1
port 5 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 10 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1363480
string GDS_START 1352726
<< end >>
