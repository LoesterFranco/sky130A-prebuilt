magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 23 380 89 649
rect 125 424 163 596
rect 125 390 127 424
rect 161 390 163 424
rect 125 364 163 390
rect 203 364 253 649
rect 293 424 359 596
rect 293 390 309 424
rect 343 390 359 424
rect 293 377 359 390
rect 23 17 89 168
rect 125 155 161 364
rect 195 276 259 330
rect 195 242 209 276
rect 243 242 259 276
rect 195 230 259 242
rect 123 76 161 155
rect 195 17 252 168
rect 293 155 339 377
rect 399 364 433 649
rect 473 424 539 596
rect 473 390 489 424
rect 523 390 539 424
rect 473 377 539 390
rect 373 276 439 330
rect 373 242 389 276
rect 423 242 439 276
rect 373 230 439 242
rect 288 76 340 155
rect 377 17 433 168
rect 473 155 533 377
rect 579 364 613 649
rect 667 424 719 596
rect 667 390 675 424
rect 709 390 719 424
rect 567 276 633 330
rect 567 242 583 276
rect 617 242 633 276
rect 567 230 633 242
rect 470 76 533 155
rect 569 17 619 168
rect 667 155 719 390
rect 759 364 793 649
rect 833 424 899 596
rect 833 390 849 424
rect 883 390 899 424
rect 833 380 899 390
rect 833 370 905 380
rect 753 276 819 330
rect 753 242 769 276
rect 803 242 819 276
rect 753 230 819 242
rect 660 76 719 155
rect 753 17 819 168
rect 853 76 905 370
rect 939 364 973 649
rect 1013 424 1079 596
rect 1013 390 1029 424
rect 1063 402 1079 424
rect 1063 390 1085 402
rect 1013 370 1085 390
rect 951 276 1017 330
rect 951 242 967 276
rect 1001 242 1017 276
rect 951 230 1017 242
rect 953 17 1017 168
rect 1051 155 1085 370
rect 1119 364 1169 649
rect 1203 424 1266 596
rect 1203 390 1219 424
rect 1253 390 1266 424
rect 1203 364 1266 390
rect 1302 364 1359 649
rect 1409 424 1458 596
rect 1409 390 1415 424
rect 1449 390 1458 424
rect 1219 352 1266 364
rect 1119 276 1185 330
rect 1119 242 1135 276
rect 1169 242 1185 276
rect 1119 230 1185 242
rect 1219 202 1268 352
rect 1309 276 1375 330
rect 1309 242 1325 276
rect 1359 242 1375 276
rect 1309 230 1375 242
rect 1051 76 1105 155
rect 1139 17 1196 168
rect 1232 157 1268 202
rect 1232 76 1277 157
rect 1311 17 1375 168
rect 1409 76 1458 390
rect 1495 364 1561 649
rect 1601 424 1635 596
rect 1601 364 1635 390
rect 1675 364 1725 649
rect 1781 424 1815 596
rect 1781 364 1815 390
rect 1855 364 1921 649
rect 1961 424 1995 596
rect 1961 364 1995 390
rect 2035 364 2101 649
rect 2141 424 2175 596
rect 2141 364 2175 390
rect 2215 364 2281 649
rect 1505 276 2183 330
rect 1505 242 1549 276
rect 1583 242 1621 276
rect 1655 242 1693 276
rect 1727 242 1765 276
rect 1799 242 1837 276
rect 1871 242 1909 276
rect 1943 242 1981 276
rect 2015 242 2053 276
rect 2087 242 2125 276
rect 2159 242 2183 276
rect 1505 230 2183 242
rect 1497 17 1965 142
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 127 390 161 424
rect 309 390 343 424
rect 209 242 243 276
rect 489 390 523 424
rect 389 242 423 276
rect 675 390 709 424
rect 583 242 617 276
rect 849 390 883 424
rect 769 242 803 276
rect 1029 390 1063 424
rect 967 242 1001 276
rect 1219 390 1253 424
rect 1415 390 1449 424
rect 1135 242 1169 276
rect 1325 242 1359 276
rect 1601 390 1635 424
rect 1781 390 1815 424
rect 1961 390 1995 424
rect 2141 390 2175 424
rect 1549 242 1583 276
rect 1621 242 1655 276
rect 1693 242 1727 276
rect 1765 242 1799 276
rect 1837 242 1871 276
rect 1909 242 1943 276
rect 1981 242 2015 276
rect 2053 242 2087 276
rect 2125 242 2159 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 115 424 2187 430
rect 115 390 127 424
rect 161 390 309 424
rect 343 390 489 424
rect 523 390 675 424
rect 709 390 849 424
rect 883 390 1029 424
rect 1063 390 1219 424
rect 1253 390 1415 424
rect 1449 390 1601 424
rect 1635 390 1781 424
rect 1815 390 1961 424
rect 1995 390 2141 424
rect 2175 390 2187 424
rect 115 384 2187 390
rect 197 276 2187 282
rect 197 242 209 276
rect 243 242 389 276
rect 423 242 583 276
rect 617 242 769 276
rect 803 242 967 276
rect 1001 242 1135 276
rect 1169 242 1325 276
rect 1359 242 1549 276
rect 1583 242 1621 276
rect 1655 242 1693 276
rect 1727 242 1765 276
rect 1799 242 1837 276
rect 1871 242 1909 276
rect 1943 242 1981 276
rect 2015 242 2053 276
rect 2087 242 2125 276
rect 2159 242 2187 276
rect 197 236 2187 242
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
rlabel metal1 s 197 236 2187 282 6 A
port 1 nsew signal input
rlabel metal1 s 115 384 2187 430 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -49 2304 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2304 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3350670
string GDS_START 3332258
<< end >>
