magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 3302 704
<< pwell >>
rect 0 0 3264 49
<< scnmos >>
rect 127 90 157 174
rect 205 90 235 174
rect 403 113 433 197
rect 503 113 533 197
rect 581 113 611 197
rect 667 113 697 197
rect 943 125 973 209
rect 1045 125 1075 209
rect 1123 125 1153 209
rect 1321 74 1351 222
rect 1519 74 1549 222
rect 1717 118 1747 202
rect 1865 118 1895 202
rect 1972 118 2002 202
rect 2136 74 2166 202
rect 2361 74 2391 202
rect 2433 74 2463 202
rect 2535 74 2565 158
rect 2613 74 2643 158
rect 2816 74 2846 202
rect 3014 78 3044 226
rect 3150 78 3180 226
<< pmoshvt >>
rect 86 464 116 592
rect 164 464 194 592
rect 390 464 420 592
rect 526 464 556 592
rect 610 464 640 592
rect 700 464 730 592
rect 915 462 945 590
rect 1038 462 1068 590
rect 1116 462 1146 590
rect 1318 368 1348 592
rect 1596 368 1626 592
rect 1801 508 1831 592
rect 1901 508 1931 592
rect 1987 508 2017 592
rect 2096 398 2126 566
rect 2315 392 2345 592
rect 2510 392 2540 592
rect 2617 508 2647 592
rect 2701 508 2731 592
rect 2843 392 2873 592
rect 3045 368 3075 592
rect 3145 368 3175 592
<< ndiff >>
rect 27 146 127 174
rect 27 112 82 146
rect 116 112 127 146
rect 27 90 127 112
rect 157 90 205 174
rect 235 149 292 174
rect 235 115 246 149
rect 280 115 292 149
rect 235 90 292 115
rect 346 172 403 197
rect 346 138 358 172
rect 392 138 403 172
rect 346 113 403 138
rect 433 172 503 197
rect 433 138 458 172
rect 492 138 503 172
rect 433 113 503 138
rect 533 113 581 197
rect 611 172 667 197
rect 611 138 622 172
rect 656 138 667 172
rect 611 113 667 138
rect 697 172 768 197
rect 697 138 722 172
rect 756 138 768 172
rect 697 113 768 138
rect 886 184 943 209
rect 886 150 898 184
rect 932 150 943 184
rect 886 125 943 150
rect 973 178 1045 209
rect 973 144 998 178
rect 1032 144 1045 178
rect 973 125 1045 144
rect 1075 125 1123 209
rect 1153 178 1210 209
rect 1153 144 1164 178
rect 1198 144 1210 178
rect 1153 125 1210 144
rect 1264 153 1321 222
rect 1264 119 1276 153
rect 1310 119 1321 153
rect 1264 74 1321 119
rect 1351 202 1408 222
rect 1351 168 1362 202
rect 1396 168 1408 202
rect 1351 120 1408 168
rect 1351 86 1362 120
rect 1396 86 1408 120
rect 1351 74 1408 86
rect 1462 127 1519 222
rect 1462 93 1474 127
rect 1508 93 1519 127
rect 1462 74 1519 93
rect 1549 210 1606 222
rect 1549 176 1560 210
rect 1594 176 1606 210
rect 1549 120 1606 176
rect 1549 86 1560 120
rect 1594 86 1606 120
rect 1660 179 1717 202
rect 1660 145 1672 179
rect 1706 145 1717 179
rect 1660 118 1717 145
rect 1747 174 1865 202
rect 1747 140 1814 174
rect 1848 140 1865 174
rect 1747 118 1865 140
rect 1895 118 1972 202
rect 2002 120 2136 202
rect 2002 118 2036 120
rect 1549 74 1606 86
rect 2017 86 2036 118
rect 2070 86 2136 120
rect 2017 74 2136 86
rect 2166 179 2226 202
rect 2166 145 2180 179
rect 2214 145 2226 179
rect 2166 74 2226 145
rect 2304 120 2361 202
rect 2304 86 2316 120
rect 2350 86 2361 120
rect 2304 74 2361 86
rect 2391 74 2433 202
rect 2463 188 2520 202
rect 2463 154 2474 188
rect 2508 158 2520 188
rect 2766 158 2816 202
rect 2508 154 2535 158
rect 2463 120 2535 154
rect 2463 86 2474 120
rect 2508 86 2535 120
rect 2463 74 2535 86
rect 2565 74 2613 158
rect 2643 120 2816 158
rect 2643 86 2654 120
rect 2688 86 2757 120
rect 2791 86 2816 120
rect 2643 74 2816 86
rect 2846 190 2903 202
rect 2846 156 2857 190
rect 2891 156 2903 190
rect 2846 120 2903 156
rect 2846 86 2857 120
rect 2891 86 2903 120
rect 2846 74 2903 86
rect 2957 191 3014 226
rect 2957 157 2969 191
rect 3003 157 3014 191
rect 2957 78 3014 157
rect 3044 214 3150 226
rect 3044 180 3105 214
rect 3139 180 3150 214
rect 3044 124 3150 180
rect 3044 90 3105 124
rect 3139 90 3150 124
rect 3044 78 3150 90
rect 3180 214 3237 226
rect 3180 180 3191 214
rect 3225 180 3237 214
rect 3180 124 3237 180
rect 3180 90 3191 124
rect 3225 90 3237 124
rect 3180 78 3237 90
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 464 86 476
rect 116 464 164 592
rect 194 578 253 592
rect 194 544 207 578
rect 241 544 253 578
rect 194 464 253 544
rect 331 520 390 592
rect 331 486 343 520
rect 377 486 390 520
rect 331 464 390 486
rect 420 580 526 592
rect 420 546 479 580
rect 513 546 526 580
rect 420 464 526 546
rect 556 464 610 592
rect 640 580 700 592
rect 640 546 653 580
rect 687 546 700 580
rect 640 512 700 546
rect 640 478 653 512
rect 687 478 700 512
rect 640 464 700 478
rect 730 580 789 592
rect 2239 596 2297 608
rect 730 546 743 580
rect 777 546 789 580
rect 730 510 789 546
rect 730 476 743 510
rect 777 476 789 510
rect 730 464 789 476
rect 843 519 915 590
rect 843 485 855 519
rect 889 485 915 519
rect 843 462 915 485
rect 945 577 1038 590
rect 945 543 991 577
rect 1025 543 1038 577
rect 945 462 1038 543
rect 1068 462 1116 590
rect 1146 578 1205 590
rect 1146 544 1159 578
rect 1193 544 1205 578
rect 1146 508 1205 544
rect 1146 474 1159 508
rect 1193 474 1205 508
rect 1146 462 1205 474
rect 1259 580 1318 592
rect 1259 546 1271 580
rect 1305 546 1318 580
rect 1259 368 1318 546
rect 1348 421 1407 592
rect 1537 580 1596 592
rect 1537 546 1549 580
rect 1583 546 1596 580
rect 1348 387 1361 421
rect 1395 387 1407 421
rect 1348 368 1407 387
rect 1537 368 1596 546
rect 1626 421 1685 592
rect 1739 580 1801 592
rect 1739 546 1752 580
rect 1786 546 1801 580
rect 1739 508 1801 546
rect 1831 567 1901 592
rect 1831 533 1854 567
rect 1888 533 1901 567
rect 1831 508 1901 533
rect 1931 508 1987 592
rect 2017 580 2078 592
rect 2017 546 2032 580
rect 2066 566 2078 580
rect 2066 546 2096 566
rect 2017 508 2096 546
rect 1626 387 1639 421
rect 1673 387 1685 421
rect 1626 368 1685 387
rect 2043 398 2096 508
rect 2126 444 2185 566
rect 2126 410 2139 444
rect 2173 410 2185 444
rect 2126 398 2185 410
rect 2239 562 2251 596
rect 2285 592 2297 596
rect 2285 562 2315 592
rect 2239 392 2315 562
rect 2345 392 2510 592
rect 2540 567 2617 592
rect 2540 533 2553 567
rect 2587 533 2617 567
rect 2540 508 2617 533
rect 2647 508 2701 592
rect 2731 580 2843 592
rect 2731 546 2770 580
rect 2804 546 2843 580
rect 2731 508 2843 546
rect 2540 392 2599 508
rect 2790 392 2843 508
rect 2873 580 2932 592
rect 2873 546 2886 580
rect 2920 546 2932 580
rect 2873 509 2932 546
rect 2873 475 2886 509
rect 2920 475 2932 509
rect 2873 438 2932 475
rect 2873 404 2886 438
rect 2920 404 2932 438
rect 2873 392 2932 404
rect 2986 580 3045 592
rect 2986 546 2998 580
rect 3032 546 3045 580
rect 2986 497 3045 546
rect 2986 463 2998 497
rect 3032 463 3045 497
rect 2986 414 3045 463
rect 2986 380 2998 414
rect 3032 380 3045 414
rect 2986 368 3045 380
rect 3075 580 3145 592
rect 3075 546 3088 580
rect 3122 546 3145 580
rect 3075 497 3145 546
rect 3075 463 3088 497
rect 3122 463 3145 497
rect 3075 414 3145 463
rect 3075 380 3088 414
rect 3122 380 3145 414
rect 3075 368 3145 380
rect 3175 580 3234 592
rect 3175 546 3188 580
rect 3222 546 3234 580
rect 3175 497 3234 546
rect 3175 463 3188 497
rect 3222 463 3234 497
rect 3175 414 3234 463
rect 3175 380 3188 414
rect 3222 380 3234 414
rect 3175 368 3234 380
<< ndiffc >>
rect 82 112 116 146
rect 246 115 280 149
rect 358 138 392 172
rect 458 138 492 172
rect 622 138 656 172
rect 722 138 756 172
rect 898 150 932 184
rect 998 144 1032 178
rect 1164 144 1198 178
rect 1276 119 1310 153
rect 1362 168 1396 202
rect 1362 86 1396 120
rect 1474 93 1508 127
rect 1560 176 1594 210
rect 1560 86 1594 120
rect 1672 145 1706 179
rect 1814 140 1848 174
rect 2036 86 2070 120
rect 2180 145 2214 179
rect 2316 86 2350 120
rect 2474 154 2508 188
rect 2474 86 2508 120
rect 2654 86 2688 120
rect 2757 86 2791 120
rect 2857 156 2891 190
rect 2857 86 2891 120
rect 2969 157 3003 191
rect 3105 180 3139 214
rect 3105 90 3139 124
rect 3191 180 3225 214
rect 3191 90 3225 124
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 207 544 241 578
rect 343 486 377 520
rect 479 546 513 580
rect 653 546 687 580
rect 653 478 687 512
rect 743 546 777 580
rect 743 476 777 510
rect 855 485 889 519
rect 991 543 1025 577
rect 1159 544 1193 578
rect 1159 474 1193 508
rect 1271 546 1305 580
rect 1549 546 1583 580
rect 1361 387 1395 421
rect 1752 546 1786 580
rect 1854 533 1888 567
rect 2032 546 2066 580
rect 1639 387 1673 421
rect 2139 410 2173 444
rect 2251 562 2285 596
rect 2553 533 2587 567
rect 2770 546 2804 580
rect 2886 546 2920 580
rect 2886 475 2920 509
rect 2886 404 2920 438
rect 2998 546 3032 580
rect 2998 463 3032 497
rect 2998 380 3032 414
rect 3088 546 3122 580
rect 3088 463 3122 497
rect 3088 380 3122 414
rect 3188 546 3222 580
rect 3188 463 3222 497
rect 3188 380 3222 414
<< poly >>
rect 86 592 116 618
rect 164 592 194 618
rect 390 592 420 618
rect 526 592 556 618
rect 610 592 640 618
rect 697 607 948 637
rect 700 592 730 607
rect 912 605 948 607
rect 915 590 945 605
rect 1038 590 1068 616
rect 1116 590 1146 616
rect 1318 592 1348 618
rect 1596 592 1626 618
rect 1801 592 1831 618
rect 1901 592 1931 618
rect 1987 592 2017 618
rect 86 449 116 464
rect 164 449 194 464
rect 390 449 420 464
rect 526 449 556 464
rect 610 449 640 464
rect 83 346 119 449
rect 161 424 197 449
rect 161 408 271 424
rect 161 394 221 408
rect 205 374 221 394
rect 255 374 271 408
rect 83 330 157 346
rect 83 296 107 330
rect 141 296 157 330
rect 83 262 157 296
rect 205 340 271 374
rect 387 419 559 449
rect 387 356 417 419
rect 607 371 643 449
rect 700 438 730 464
rect 915 447 945 462
rect 1038 447 1068 462
rect 1116 447 1146 462
rect 205 306 221 340
rect 255 306 271 340
rect 205 290 271 306
rect 351 340 417 356
rect 351 306 367 340
rect 401 306 417 340
rect 351 290 417 306
rect 467 355 533 371
rect 467 321 483 355
rect 517 321 533 355
rect 467 305 533 321
rect 575 355 643 371
rect 575 321 591 355
rect 625 321 643 355
rect 575 305 643 321
rect 798 404 864 420
rect 798 370 814 404
rect 848 370 864 404
rect 798 336 864 370
rect 912 356 948 447
rect 83 228 107 262
rect 141 228 157 262
rect 351 242 381 290
rect 83 212 157 228
rect 127 174 157 212
rect 205 212 433 242
rect 205 174 235 212
rect 403 197 433 212
rect 503 197 533 305
rect 581 197 611 305
rect 798 302 814 336
rect 848 302 864 336
rect 798 268 864 302
rect 907 340 973 356
rect 907 306 923 340
rect 957 306 973 340
rect 907 290 973 306
rect 1035 302 1071 447
rect 1113 424 1149 447
rect 1113 408 1179 424
rect 1113 374 1129 408
rect 1163 374 1179 408
rect 1113 358 1179 374
rect 1439 412 1505 428
rect 1439 378 1455 412
rect 1489 378 1505 412
rect 1318 353 1348 368
rect 1439 353 1505 378
rect 2096 566 2126 592
rect 1801 493 1831 508
rect 1901 493 1931 508
rect 1987 493 2017 508
rect 1798 476 1834 493
rect 1717 460 1834 476
rect 1717 426 1733 460
rect 1767 446 1834 460
rect 1898 451 1934 493
rect 1767 426 1783 446
rect 1717 410 1783 426
rect 1876 435 1942 451
rect 1876 401 1892 435
rect 1926 401 1942 435
rect 1876 385 1942 401
rect 1876 368 1906 385
rect 1596 353 1626 368
rect 1717 353 1906 368
rect 1315 310 1351 353
rect 1439 338 1906 353
rect 1439 323 1747 338
rect 798 242 814 268
rect 667 234 814 242
rect 848 234 864 268
rect 667 212 864 234
rect 667 197 697 212
rect 798 200 864 212
rect 943 209 973 290
rect 1015 286 1081 302
rect 1015 252 1031 286
rect 1065 252 1081 286
rect 1015 236 1081 252
rect 1315 294 1381 310
rect 1315 260 1331 294
rect 1365 260 1381 294
rect 1315 244 1381 260
rect 1045 209 1075 236
rect 1123 209 1153 235
rect 1321 222 1351 244
rect 1519 222 1549 323
rect 798 166 814 200
rect 848 166 864 200
rect 798 132 864 166
rect 127 64 157 90
rect 205 64 235 90
rect 403 87 433 113
rect 503 87 533 113
rect 581 87 611 113
rect 667 87 697 113
rect 798 98 814 132
rect 848 98 864 132
rect 798 82 864 98
rect 943 51 973 125
rect 1045 99 1075 125
rect 1123 51 1153 125
rect 1717 202 1747 323
rect 1984 297 2020 493
rect 2315 592 2345 618
rect 2510 592 2540 618
rect 2617 592 2647 618
rect 2701 592 2731 618
rect 2843 592 2873 618
rect 3045 592 3075 618
rect 3145 592 3175 618
rect 2096 383 2126 398
rect 2617 493 2647 508
rect 2701 493 2731 508
rect 2614 408 2650 493
rect 2698 476 2734 493
rect 2692 460 2758 476
rect 2692 426 2708 460
rect 2742 426 2758 460
rect 2692 410 2758 426
rect 2093 366 2129 383
rect 2315 377 2345 392
rect 2510 377 2540 392
rect 2080 350 2166 366
rect 2080 316 2096 350
rect 2130 316 2166 350
rect 2080 300 2166 316
rect 2312 304 2348 377
rect 2507 360 2543 377
rect 1864 274 1930 290
rect 1864 240 1880 274
rect 1914 240 1930 274
rect 1864 224 1930 240
rect 1972 281 2038 297
rect 1972 247 1988 281
rect 2022 247 2038 281
rect 1972 231 2038 247
rect 1865 202 1895 224
rect 1972 202 2002 231
rect 2136 202 2166 300
rect 2214 288 2348 304
rect 2390 344 2463 360
rect 2390 310 2406 344
rect 2440 310 2463 344
rect 2390 294 2463 310
rect 2505 344 2571 360
rect 2505 310 2521 344
rect 2555 310 2571 344
rect 2620 311 2650 408
rect 2505 294 2571 310
rect 2613 295 2679 311
rect 2214 254 2230 288
rect 2264 254 2298 288
rect 2332 254 2348 288
rect 2214 252 2348 254
rect 2214 222 2391 252
rect 2361 202 2391 222
rect 2433 202 2463 294
rect 1717 92 1747 118
rect 1865 92 1895 118
rect 1972 92 2002 118
rect 2535 158 2565 294
rect 2613 261 2629 295
rect 2663 261 2679 295
rect 2613 245 2679 261
rect 2721 203 2751 410
rect 2843 377 2873 392
rect 2840 306 2876 377
rect 3045 353 3075 368
rect 3145 353 3175 368
rect 2793 290 2876 306
rect 2793 256 2809 290
rect 2843 271 2876 290
rect 3042 271 3078 353
rect 3142 330 3178 353
rect 2843 256 3078 271
rect 3120 314 3186 330
rect 3120 280 3136 314
rect 3170 280 3186 314
rect 3120 264 3186 280
rect 2793 241 3078 256
rect 2793 240 2870 241
rect 2613 173 2751 203
rect 2816 202 2846 240
rect 3014 226 3044 241
rect 3150 226 3180 264
rect 2613 158 2643 173
rect 943 21 1153 51
rect 1321 48 1351 74
rect 1519 48 1549 74
rect 2136 48 2166 74
rect 2361 48 2391 74
rect 2433 48 2463 74
rect 2535 48 2565 74
rect 2613 48 2643 74
rect 2816 48 2846 74
rect 3014 52 3044 78
rect 3150 52 3180 78
<< polycont >>
rect 221 374 255 408
rect 107 296 141 330
rect 221 306 255 340
rect 367 306 401 340
rect 483 321 517 355
rect 591 321 625 355
rect 814 370 848 404
rect 107 228 141 262
rect 814 302 848 336
rect 923 306 957 340
rect 1129 374 1163 408
rect 1455 378 1489 412
rect 1733 426 1767 460
rect 1892 401 1926 435
rect 814 234 848 268
rect 1031 252 1065 286
rect 1331 260 1365 294
rect 814 166 848 200
rect 814 98 848 132
rect 2708 426 2742 460
rect 2096 316 2130 350
rect 1880 240 1914 274
rect 1988 247 2022 281
rect 2406 310 2440 344
rect 2521 310 2555 344
rect 2230 254 2264 288
rect 2298 254 2332 288
rect 2629 261 2663 295
rect 2809 256 2843 290
rect 3136 280 3170 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 191 578 241 649
rect 191 544 207 578
rect 191 526 241 544
rect 275 581 445 615
rect 23 476 39 510
rect 73 492 89 510
rect 275 492 309 581
rect 73 476 309 492
rect 23 458 309 476
rect 343 520 377 547
rect 23 162 57 458
rect 343 424 377 486
rect 411 496 445 581
rect 479 580 529 649
rect 513 546 529 580
rect 479 530 529 546
rect 637 580 709 596
rect 637 546 653 580
rect 687 546 709 580
rect 637 512 709 546
rect 637 496 653 512
rect 411 478 653 496
rect 687 478 709 512
rect 411 462 709 478
rect 575 424 641 428
rect 205 408 533 424
rect 205 374 221 408
rect 255 390 533 408
rect 255 374 271 390
rect 91 330 167 356
rect 91 296 107 330
rect 141 296 167 330
rect 91 262 167 296
rect 91 228 107 262
rect 141 228 167 262
rect 91 212 167 228
rect 205 340 271 374
rect 205 306 221 340
rect 255 306 271 340
rect 205 256 271 306
rect 313 340 417 356
rect 313 306 367 340
rect 401 306 417 340
rect 313 290 417 306
rect 467 355 533 390
rect 467 321 483 355
rect 517 321 533 355
rect 467 305 533 321
rect 575 390 607 424
rect 575 355 641 390
rect 575 321 591 355
rect 625 321 641 355
rect 575 305 641 321
rect 675 269 709 462
rect 205 222 408 256
rect 23 146 132 162
rect 23 112 82 146
rect 116 112 132 146
rect 23 96 132 112
rect 230 149 296 178
rect 230 115 246 149
rect 280 115 296 149
rect 230 17 296 115
rect 342 172 408 222
rect 606 235 709 269
rect 743 581 957 615
rect 743 580 793 581
rect 777 546 793 580
rect 743 510 793 546
rect 777 476 793 510
rect 743 460 793 476
rect 827 519 889 547
rect 827 485 855 519
rect 342 138 358 172
rect 392 138 408 172
rect 342 109 408 138
rect 442 172 508 201
rect 442 138 458 172
rect 492 138 508 172
rect 442 17 508 138
rect 606 172 672 235
rect 743 201 777 460
rect 827 458 889 485
rect 923 492 957 581
rect 991 577 1041 649
rect 1025 543 1041 577
rect 991 526 1041 543
rect 1143 578 1209 594
rect 1143 544 1159 578
rect 1193 544 1209 578
rect 1143 508 1209 544
rect 1255 580 1321 649
rect 1255 546 1271 580
rect 1305 546 1321 580
rect 1255 530 1321 546
rect 1533 580 1599 649
rect 1533 546 1549 580
rect 1583 546 1599 580
rect 1533 530 1599 546
rect 1633 580 1804 596
rect 1633 546 1752 580
rect 1786 546 1804 580
rect 1838 567 1904 596
rect 1143 492 1159 508
rect 923 474 1159 492
rect 1193 496 1209 508
rect 1633 496 1667 546
rect 1838 533 1854 567
rect 1888 533 1904 567
rect 2016 580 2082 649
rect 2016 546 2032 580
rect 2066 546 2082 580
rect 2235 596 2301 649
rect 2235 562 2251 596
rect 2285 562 2301 596
rect 2235 546 2301 562
rect 2553 567 2639 596
rect 1838 512 1904 533
rect 2587 533 2639 567
rect 1193 474 1667 496
rect 1808 478 1904 512
rect 1938 478 2519 512
rect 2553 504 2639 533
rect 2728 580 2846 649
rect 2728 546 2770 580
rect 2804 546 2846 580
rect 2728 530 2846 546
rect 2886 580 2920 596
rect 923 462 1667 474
rect 923 458 1242 462
rect 827 424 861 458
rect 606 138 622 172
rect 656 138 672 172
rect 606 109 672 138
rect 706 172 777 201
rect 706 138 722 172
rect 756 138 777 172
rect 706 109 777 138
rect 811 408 1174 424
rect 811 404 1129 408
rect 811 370 814 404
rect 848 390 1129 404
rect 848 370 861 390
rect 811 336 861 370
rect 1113 374 1129 390
rect 1163 374 1174 408
rect 1113 358 1174 374
rect 811 302 814 336
rect 848 302 861 336
rect 811 268 861 302
rect 895 340 973 356
rect 895 306 923 340
rect 957 306 973 340
rect 895 290 973 306
rect 811 234 814 268
rect 848 234 861 268
rect 1015 286 1127 302
rect 1015 252 1031 286
rect 1065 252 1127 286
rect 1015 236 1127 252
rect 811 213 861 234
rect 811 200 948 213
rect 1208 202 1242 458
rect 1345 421 1505 428
rect 1345 387 1361 421
rect 1395 412 1505 421
rect 1395 387 1455 412
rect 1345 378 1455 387
rect 1489 378 1505 412
rect 1345 364 1505 378
rect 1411 362 1505 364
rect 1315 294 1415 310
rect 1315 260 1331 294
rect 1365 260 1415 294
rect 1315 236 1415 260
rect 1471 202 1505 362
rect 1555 330 1589 462
rect 1717 460 1774 476
rect 1717 428 1733 460
rect 1623 426 1733 428
rect 1767 426 1774 460
rect 1623 421 1774 426
rect 1623 387 1639 421
rect 1673 387 1774 421
rect 1623 364 1774 387
rect 1555 296 1706 330
rect 811 166 814 200
rect 848 184 948 200
rect 848 166 898 184
rect 811 150 898 166
rect 932 150 948 184
rect 811 132 948 150
rect 811 98 814 132
rect 848 121 948 132
rect 982 178 1048 202
rect 982 144 998 178
rect 1032 144 1048 178
rect 848 98 861 121
rect 811 82 861 98
rect 982 17 1048 144
rect 1148 178 1242 202
rect 1148 144 1164 178
rect 1198 144 1242 178
rect 1148 121 1242 144
rect 1276 153 1310 202
rect 1276 17 1310 119
rect 1346 168 1362 202
rect 1396 168 1505 202
rect 1560 210 1610 226
rect 1594 176 1610 210
rect 1346 120 1412 168
rect 1346 86 1362 120
rect 1396 86 1412 120
rect 1346 70 1412 86
rect 1458 127 1524 134
rect 1458 93 1474 127
rect 1508 93 1524 127
rect 1458 17 1524 93
rect 1560 120 1610 176
rect 1594 86 1610 120
rect 1656 179 1706 296
rect 1656 145 1672 179
rect 1656 119 1706 145
rect 1560 85 1610 86
rect 1740 85 1774 364
rect 1808 358 1842 478
rect 1938 444 1972 478
rect 1876 435 1972 444
rect 1876 401 1892 435
rect 1926 401 1972 435
rect 2123 410 2139 444
rect 2173 410 2214 444
rect 1876 392 1972 401
rect 2080 358 2146 366
rect 1808 350 2146 358
rect 1808 324 2096 350
rect 1808 190 1842 324
rect 2080 316 2096 324
rect 2130 316 2146 350
rect 2080 306 2146 316
rect 2180 304 2214 410
rect 2485 360 2519 478
rect 2605 377 2639 504
rect 2886 509 2920 546
rect 2692 475 2886 476
rect 2692 460 2920 475
rect 2692 426 2708 460
rect 2742 438 2920 460
rect 2742 426 2886 438
rect 2692 424 2886 426
rect 2692 411 2815 424
rect 2809 390 2815 411
rect 2849 404 2886 424
rect 2849 390 2920 404
rect 2809 384 2920 390
rect 2390 344 2451 360
rect 2390 310 2406 344
rect 2440 310 2451 344
rect 1876 274 1938 290
rect 1876 240 1880 274
rect 1914 240 1938 274
rect 1876 224 1938 240
rect 1972 281 2038 290
rect 1972 247 1988 281
rect 2022 272 2038 281
rect 2180 288 2348 304
rect 2180 272 2230 288
rect 2022 254 2230 272
rect 2264 254 2298 288
rect 2332 254 2348 288
rect 2022 247 2348 254
rect 1972 238 2348 247
rect 2390 260 2451 310
rect 2485 344 2571 360
rect 2485 310 2521 344
rect 2555 310 2571 344
rect 2605 343 2775 377
rect 2485 294 2571 310
rect 2613 295 2679 309
rect 2613 261 2629 295
rect 2663 261 2679 295
rect 2613 260 2679 261
rect 1898 204 1938 224
rect 1808 174 1864 190
rect 1808 140 1814 174
rect 1848 140 1864 174
rect 1808 124 1864 140
rect 1898 170 2146 204
rect 1898 85 1938 170
rect 1560 51 1938 85
rect 2013 120 2078 136
rect 2013 86 2036 120
rect 2070 86 2078 120
rect 2013 17 2078 86
rect 2112 85 2146 170
rect 2180 179 2214 238
rect 2390 226 2679 260
rect 2741 306 2775 343
rect 2741 290 2852 306
rect 2741 256 2809 290
rect 2843 256 2852 290
rect 2741 240 2852 256
rect 2390 204 2424 226
rect 2180 119 2214 145
rect 2248 170 2424 204
rect 2741 188 2775 240
rect 2886 206 2920 384
rect 2248 85 2282 170
rect 2458 154 2474 188
rect 2508 154 2775 188
rect 2841 190 2920 206
rect 2841 156 2857 190
rect 2891 156 2920 190
rect 2112 51 2282 85
rect 2316 120 2366 136
rect 2350 86 2366 120
rect 2316 17 2366 86
rect 2458 120 2524 154
rect 2841 120 2920 156
rect 2969 580 3048 596
rect 2969 546 2998 580
rect 3032 546 3048 580
rect 2969 497 3048 546
rect 2969 463 2998 497
rect 3032 463 3048 497
rect 2969 414 3048 463
rect 2969 380 2998 414
rect 3032 380 3048 414
rect 2969 364 3048 380
rect 3088 580 3138 649
rect 3122 546 3138 580
rect 3088 497 3138 546
rect 3122 463 3138 497
rect 3088 414 3138 463
rect 3122 380 3138 414
rect 3088 364 3138 380
rect 3172 580 3247 596
rect 3172 546 3188 580
rect 3222 546 3247 580
rect 3172 497 3247 546
rect 3172 463 3188 497
rect 3222 463 3247 497
rect 3172 414 3247 463
rect 3172 380 3188 414
rect 3222 380 3247 414
rect 3172 364 3247 380
rect 2969 191 3003 364
rect 2969 124 3003 157
rect 3037 314 3179 330
rect 3037 280 3136 314
rect 3170 280 3179 314
rect 3037 264 3179 280
rect 2458 86 2474 120
rect 2508 86 2524 120
rect 2458 70 2524 86
rect 2638 86 2654 120
rect 2688 86 2757 120
rect 2791 86 2807 120
rect 2638 17 2807 86
rect 2841 86 2857 120
rect 2891 86 2920 120
rect 2841 85 2920 86
rect 3037 85 3071 264
rect 3213 230 3247 364
rect 2841 51 3071 85
rect 3105 214 3139 230
rect 3105 124 3139 180
rect 3105 17 3139 90
rect 3175 214 3247 230
rect 3175 180 3191 214
rect 3225 180 3247 214
rect 3175 124 3247 180
rect 3175 90 3191 124
rect 3225 90 3247 124
rect 3175 74 3247 90
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 607 390 641 424
rect 2815 390 2849 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
<< metal1 >>
rect 0 683 3264 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 0 617 3264 649
rect 595 424 653 430
rect 595 390 607 424
rect 641 421 653 424
rect 2803 424 2861 430
rect 2803 421 2815 424
rect 641 393 2815 421
rect 641 390 653 393
rect 595 384 653 390
rect 2803 390 2815 393
rect 2849 390 2861 424
rect 2803 384 2861 390
rect 0 17 3264 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
rect 0 -49 3264 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sedfxbp_1
flabel comment s 1657 341 1657 341 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 3264 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 3264 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 0 617 3264 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 3264 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 3199 390 3233 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 3199 464 3233 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 3199 538 3233 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 3007 390 3041 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3007 464 3041 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 3007 538 3041 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 1087 242 1121 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 DE
port 3 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 3264 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 476332
string GDS_START 453500
<< end >>
