magic
tech sky130A
magscale 1 2
timestamp 1599588209
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 0 0 1152 49
<< scpmos >>
rect 86 387 116 587
rect 186 387 216 587
rect 276 387 306 587
rect 376 387 406 587
rect 484 387 514 555
rect 590 387 620 555
rect 736 368 766 592
rect 826 368 856 592
rect 936 368 966 592
rect 1026 368 1056 592
<< nmoslvt >>
rect 84 125 114 253
rect 185 125 215 253
rect 271 125 301 253
rect 387 125 417 253
rect 473 125 503 253
rect 559 125 589 253
rect 773 74 803 222
rect 859 74 889 222
rect 952 74 982 222
rect 1038 74 1068 222
<< ndiff >>
rect 27 241 84 253
rect 27 207 39 241
rect 73 207 84 241
rect 27 171 84 207
rect 27 137 39 171
rect 73 137 84 171
rect 27 125 84 137
rect 114 171 185 253
rect 114 137 139 171
rect 173 137 185 171
rect 114 125 185 137
rect 215 239 271 253
rect 215 205 226 239
rect 260 205 271 239
rect 215 171 271 205
rect 215 137 226 171
rect 260 137 271 171
rect 215 125 271 137
rect 301 171 387 253
rect 301 137 328 171
rect 362 137 387 171
rect 301 125 387 137
rect 417 239 473 253
rect 417 205 428 239
rect 462 205 473 239
rect 417 171 473 205
rect 417 137 428 171
rect 462 137 473 171
rect 417 125 473 137
rect 503 241 559 253
rect 503 207 514 241
rect 548 207 559 241
rect 503 171 559 207
rect 503 137 514 171
rect 548 137 559 171
rect 503 125 559 137
rect 589 178 662 253
rect 589 144 616 178
rect 650 144 662 178
rect 589 125 662 144
rect 716 185 773 222
rect 716 151 728 185
rect 762 151 773 185
rect 716 117 773 151
rect 716 83 728 117
rect 762 83 773 117
rect 716 74 773 83
rect 803 201 859 222
rect 803 167 814 201
rect 848 167 859 201
rect 803 116 859 167
rect 803 82 814 116
rect 848 82 859 116
rect 803 74 859 82
rect 889 117 952 222
rect 889 83 903 117
rect 937 83 952 117
rect 889 74 952 83
rect 982 210 1038 222
rect 982 176 993 210
rect 1027 176 1038 210
rect 982 120 1038 176
rect 982 86 993 120
rect 1027 86 1038 120
rect 982 74 1038 86
rect 1068 210 1125 222
rect 1068 176 1079 210
rect 1113 176 1125 210
rect 1068 120 1125 176
rect 1068 86 1079 120
rect 1113 86 1125 120
rect 1068 74 1125 86
<< pdiff >>
rect 27 575 86 587
rect 27 541 39 575
rect 73 541 86 575
rect 27 504 86 541
rect 27 470 39 504
rect 73 470 86 504
rect 27 433 86 470
rect 27 399 39 433
rect 73 399 86 433
rect 27 387 86 399
rect 116 576 186 587
rect 116 542 139 576
rect 173 542 186 576
rect 116 508 186 542
rect 116 474 139 508
rect 173 474 186 508
rect 116 440 186 474
rect 116 406 139 440
rect 173 406 186 440
rect 116 387 186 406
rect 216 531 276 587
rect 216 497 229 531
rect 263 497 276 531
rect 216 440 276 497
rect 216 406 229 440
rect 263 406 276 440
rect 216 387 276 406
rect 306 579 376 587
rect 306 545 329 579
rect 363 545 376 579
rect 306 492 376 545
rect 306 458 329 492
rect 363 458 376 492
rect 306 387 376 458
rect 406 555 459 587
rect 683 555 736 592
rect 406 508 484 555
rect 406 474 429 508
rect 463 474 484 508
rect 406 387 484 474
rect 514 543 590 555
rect 514 509 529 543
rect 563 509 590 543
rect 514 440 590 509
rect 514 406 529 440
rect 563 406 590 440
rect 514 387 590 406
rect 620 510 736 555
rect 620 476 655 510
rect 689 476 736 510
rect 620 387 736 476
rect 683 368 736 387
rect 766 580 826 592
rect 766 546 779 580
rect 813 546 826 580
rect 766 497 826 546
rect 766 463 779 497
rect 813 463 826 497
rect 766 414 826 463
rect 766 380 779 414
rect 813 380 826 414
rect 766 368 826 380
rect 856 582 936 592
rect 856 548 879 582
rect 913 548 936 582
rect 856 514 936 548
rect 856 480 879 514
rect 913 480 936 514
rect 856 446 936 480
rect 856 412 879 446
rect 913 412 936 446
rect 856 368 936 412
rect 966 580 1026 592
rect 966 546 979 580
rect 1013 546 1026 580
rect 966 497 1026 546
rect 966 463 979 497
rect 1013 463 1026 497
rect 966 414 1026 463
rect 966 380 979 414
rect 1013 380 1026 414
rect 966 368 1026 380
rect 1056 580 1125 592
rect 1056 546 1079 580
rect 1113 546 1125 580
rect 1056 510 1125 546
rect 1056 476 1079 510
rect 1113 476 1125 510
rect 1056 440 1125 476
rect 1056 406 1079 440
rect 1113 406 1125 440
rect 1056 368 1125 406
<< ndiffc >>
rect 39 207 73 241
rect 39 137 73 171
rect 139 137 173 171
rect 226 205 260 239
rect 226 137 260 171
rect 328 137 362 171
rect 428 205 462 239
rect 428 137 462 171
rect 514 207 548 241
rect 514 137 548 171
rect 616 144 650 178
rect 728 151 762 185
rect 728 83 762 117
rect 814 167 848 201
rect 814 82 848 116
rect 903 83 937 117
rect 993 176 1027 210
rect 993 86 1027 120
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 39 541 73 575
rect 39 470 73 504
rect 39 399 73 433
rect 139 542 173 576
rect 139 474 173 508
rect 139 406 173 440
rect 229 497 263 531
rect 229 406 263 440
rect 329 545 363 579
rect 329 458 363 492
rect 429 474 463 508
rect 529 509 563 543
rect 529 406 563 440
rect 655 476 689 510
rect 779 546 813 580
rect 779 463 813 497
rect 779 380 813 414
rect 879 548 913 582
rect 879 480 913 514
rect 879 412 913 446
rect 979 546 1013 580
rect 979 463 1013 497
rect 979 380 1013 414
rect 1079 546 1113 580
rect 1079 476 1113 510
rect 1079 406 1113 440
<< poly >>
rect 86 587 116 613
rect 186 587 216 613
rect 276 587 306 613
rect 376 587 406 613
rect 736 592 766 618
rect 826 592 856 618
rect 936 592 966 618
rect 1026 592 1056 618
rect 484 555 514 581
rect 590 555 620 581
rect 86 372 116 387
rect 186 372 216 387
rect 276 372 306 387
rect 376 372 406 387
rect 484 372 514 387
rect 590 372 620 387
rect 83 268 119 372
rect 183 355 219 372
rect 273 355 309 372
rect 373 355 409 372
rect 481 355 517 372
rect 587 355 623 372
rect 167 339 309 355
rect 167 305 183 339
rect 217 305 251 339
rect 285 305 309 339
rect 167 289 309 305
rect 359 339 425 355
rect 359 305 375 339
rect 409 305 425 339
rect 359 289 425 305
rect 473 339 623 355
rect 736 353 766 368
rect 826 353 856 368
rect 936 353 966 368
rect 1026 353 1056 368
rect 473 305 505 339
rect 539 305 573 339
rect 607 305 623 339
rect 733 310 769 353
rect 823 310 859 353
rect 933 352 969 353
rect 1023 352 1059 353
rect 933 310 1059 352
rect 473 289 623 305
rect 689 294 1059 310
rect 84 253 114 268
rect 185 253 215 289
rect 271 253 301 289
rect 387 253 417 289
rect 473 253 503 289
rect 559 253 589 289
rect 689 260 705 294
rect 739 260 773 294
rect 807 260 841 294
rect 875 260 909 294
rect 943 274 1059 294
rect 943 260 1068 274
rect 689 244 1068 260
rect 773 222 803 244
rect 859 222 889 244
rect 952 222 982 244
rect 1038 222 1068 244
rect 84 51 114 125
rect 185 99 215 125
rect 271 99 301 125
rect 387 51 417 125
rect 473 99 503 125
rect 559 99 589 125
rect 84 21 417 51
rect 773 48 803 74
rect 859 48 889 74
rect 952 48 982 74
rect 1038 48 1068 74
<< polycont >>
rect 183 305 217 339
rect 251 305 285 339
rect 375 305 409 339
rect 505 305 539 339
rect 573 305 607 339
rect 705 260 739 294
rect 773 260 807 294
rect 841 260 875 294
rect 909 260 943 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 575 89 649
rect 23 541 39 575
rect 73 541 89 575
rect 23 504 89 541
rect 23 470 39 504
rect 73 470 89 504
rect 23 433 89 470
rect 23 399 39 433
rect 73 399 89 433
rect 23 383 89 399
rect 123 581 379 615
rect 123 576 173 581
rect 123 542 139 576
rect 313 579 379 581
rect 123 508 173 542
rect 123 474 139 508
rect 123 440 173 474
rect 123 406 139 440
rect 123 390 173 406
rect 213 531 279 547
rect 213 497 229 531
rect 263 497 279 531
rect 213 440 279 497
rect 313 545 329 579
rect 363 545 379 579
rect 313 492 379 545
rect 313 458 329 492
rect 363 458 379 492
rect 413 508 479 649
rect 413 474 429 508
rect 463 474 479 508
rect 413 458 479 474
rect 513 543 579 559
rect 513 509 529 543
rect 563 509 579 543
rect 213 406 229 440
rect 263 424 279 440
rect 513 440 579 509
rect 627 510 723 649
rect 627 476 655 510
rect 689 476 723 510
rect 627 460 723 476
rect 763 580 829 596
rect 763 546 779 580
rect 813 546 829 580
rect 763 497 829 546
rect 763 463 779 497
rect 813 463 829 497
rect 513 424 529 440
rect 263 406 529 424
rect 563 424 579 440
rect 563 406 715 424
rect 213 390 715 406
rect 167 339 301 356
rect 167 305 183 339
rect 217 305 251 339
rect 285 305 301 339
rect 167 289 301 305
rect 359 339 455 356
rect 359 305 375 339
rect 409 305 455 339
rect 359 289 455 305
rect 489 339 647 356
rect 489 305 505 339
rect 539 305 573 339
rect 607 305 647 339
rect 489 303 647 305
rect 681 310 715 390
rect 763 414 829 463
rect 763 380 779 414
rect 813 380 829 414
rect 863 582 929 649
rect 863 548 879 582
rect 913 548 929 582
rect 863 514 929 548
rect 863 480 879 514
rect 913 480 929 514
rect 863 446 929 480
rect 863 412 879 446
rect 913 412 929 446
rect 963 580 1029 596
rect 963 546 979 580
rect 1013 546 1029 580
rect 963 497 1029 546
rect 963 463 979 497
rect 1013 463 1029 497
rect 963 414 1029 463
rect 763 378 829 380
rect 963 380 979 414
rect 1013 380 1029 414
rect 1063 580 1129 649
rect 1063 546 1079 580
rect 1113 546 1129 580
rect 1063 510 1129 546
rect 1063 476 1079 510
rect 1113 476 1129 510
rect 1063 440 1129 476
rect 1063 406 1079 440
rect 1113 406 1129 440
rect 1063 390 1129 406
rect 963 378 1029 380
rect 763 356 1029 378
rect 763 344 1127 356
rect 993 310 1127 344
rect 681 294 959 310
rect 681 269 705 294
rect 514 260 705 269
rect 739 260 773 294
rect 807 260 841 294
rect 875 260 909 294
rect 943 260 959 294
rect 23 255 89 257
rect 23 241 478 255
rect 23 207 39 241
rect 73 239 478 241
rect 73 221 226 239
rect 73 207 89 221
rect 23 171 89 207
rect 260 221 428 239
rect 260 205 276 221
rect 23 137 39 171
rect 73 137 89 171
rect 23 121 89 137
rect 123 171 190 187
rect 123 137 139 171
rect 173 137 190 171
rect 123 17 190 137
rect 226 171 276 205
rect 412 205 428 221
rect 462 205 478 239
rect 260 137 276 171
rect 226 121 276 137
rect 312 171 378 187
rect 312 137 328 171
rect 362 137 378 171
rect 312 17 378 137
rect 412 171 478 205
rect 412 137 428 171
rect 462 137 478 171
rect 412 87 478 137
rect 514 241 959 260
rect 548 235 959 241
rect 548 207 564 235
rect 514 171 564 207
rect 993 210 1027 310
rect 548 137 564 171
rect 514 121 564 137
rect 600 178 666 201
rect 600 144 616 178
rect 650 144 666 178
rect 600 87 666 144
rect 412 53 666 87
rect 712 185 762 201
rect 712 151 728 185
rect 712 117 762 151
rect 712 83 728 117
rect 712 17 762 83
rect 798 167 814 201
rect 848 176 993 201
rect 848 167 1027 176
rect 798 116 848 167
rect 798 82 814 116
rect 798 66 848 82
rect 884 117 957 133
rect 884 83 903 117
rect 937 83 957 117
rect 884 17 957 83
rect 993 120 1027 167
rect 993 70 1027 86
rect 1063 210 1129 226
rect 1063 176 1079 210
rect 1113 176 1129 210
rect 1063 120 1129 176
rect 1063 86 1079 120
rect 1113 86 1129 120
rect 1063 17 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21a_4
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1053078
string GDS_START 1043364
<< end >>
