magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 130 582
<< psubdiff >>
rect 29 145 63 169
rect 29 64 63 111
<< nsubdiff >>
rect 29 447 63 480
rect 29 363 63 413
rect 29 305 63 329
<< psubdiffcont >>
rect 29 111 63 145
<< nsubdiffcont >>
rect 29 413 63 447
rect 29 329 63 363
<< locali >>
rect 0 527 29 561
rect 63 527 92 561
rect 17 459 75 491
rect 17 413 29 459
rect 63 413 75 459
rect 17 363 75 413
rect 17 329 29 363
rect 63 329 75 363
rect 17 294 75 329
rect 17 145 75 162
rect 17 111 29 145
rect 63 111 75 145
rect 17 17 75 111
rect 0 -17 29 17
rect 63 -17 92 17
<< viali >>
rect 29 527 63 561
rect 29 447 63 459
rect 29 425 63 447
rect 29 -17 63 17
<< metal1 >>
rect 0 561 92 592
rect 0 527 29 561
rect 63 527 92 561
rect 0 496 92 527
rect 17 459 75 465
rect 17 425 29 459
rect 63 425 75 459
rect 17 419 75 425
rect 0 17 92 48
rect 0 -17 29 17
rect 63 -17 92 17
rect 0 -48 92 -17
<< labels >>
flabel corelocali s 34 361 63 388 0 FreeSans 250 0 0 0 VPB
port 2 nsew
flabel metal1 s 32 -13 62 14 0 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel metal1 s 31 528 61 559 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
rlabel comment s 0 0 0 0 4 tapvgnd_1
<< properties >>
string FIXED_BBOX 0 0 92 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 953976
string GDS_START 952104
string path 0.000 0.000 2.300 0.000 
<< end >>
