magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 127 368 163 568
rect 211 368 247 568
rect 325 368 361 568
rect 463 368 499 592
rect 553 368 589 592
<< nmoslvt >>
rect 125 74 155 222
rect 247 74 277 222
rect 342 74 372 222
rect 568 74 598 222
rect 654 74 684 222
<< ndiff >>
rect 54 202 125 222
rect 54 168 66 202
rect 100 168 125 202
rect 54 118 125 168
rect 54 84 66 118
rect 100 84 125 118
rect 54 74 125 84
rect 155 120 247 222
rect 155 86 181 120
rect 215 86 247 120
rect 155 74 247 86
rect 277 202 342 222
rect 277 168 297 202
rect 331 168 342 202
rect 277 118 342 168
rect 277 84 297 118
rect 331 84 342 118
rect 277 74 342 84
rect 372 186 443 222
rect 372 152 383 186
rect 417 152 443 186
rect 372 118 443 152
rect 372 84 383 118
rect 417 84 443 118
rect 372 74 443 84
rect 497 194 568 222
rect 497 160 509 194
rect 543 160 568 194
rect 497 120 568 160
rect 497 86 509 120
rect 543 86 568 120
rect 497 74 568 86
rect 598 210 654 222
rect 598 176 609 210
rect 643 176 654 210
rect 598 120 654 176
rect 598 86 609 120
rect 643 86 654 120
rect 598 74 654 86
rect 684 210 741 222
rect 684 176 695 210
rect 729 176 741 210
rect 684 120 741 176
rect 684 86 695 120
rect 729 86 741 120
rect 684 74 741 86
<< pdiff >>
rect 389 582 463 592
rect 389 568 409 582
rect 71 556 127 568
rect 71 522 83 556
rect 117 522 127 556
rect 71 485 127 522
rect 71 451 83 485
rect 117 451 127 485
rect 71 414 127 451
rect 71 380 83 414
rect 117 380 127 414
rect 71 368 127 380
rect 163 368 211 568
rect 247 556 325 568
rect 247 522 281 556
rect 315 522 325 556
rect 247 485 325 522
rect 247 451 281 485
rect 315 451 325 485
rect 247 414 325 451
rect 247 380 281 414
rect 315 380 325 414
rect 247 368 325 380
rect 361 548 409 568
rect 443 548 463 582
rect 361 514 463 548
rect 361 480 409 514
rect 443 480 463 514
rect 361 446 463 480
rect 361 412 409 446
rect 443 412 463 446
rect 361 368 463 412
rect 499 580 553 592
rect 499 546 509 580
rect 543 546 553 580
rect 499 497 553 546
rect 499 463 509 497
rect 543 463 553 497
rect 499 414 553 463
rect 499 380 509 414
rect 543 380 553 414
rect 499 368 553 380
rect 589 580 655 592
rect 589 546 609 580
rect 643 546 655 580
rect 589 462 655 546
rect 589 428 609 462
rect 643 428 655 462
rect 589 368 655 428
<< ndiffc >>
rect 66 168 100 202
rect 66 84 100 118
rect 181 86 215 120
rect 297 168 331 202
rect 297 84 331 118
rect 383 152 417 186
rect 383 84 417 118
rect 509 160 543 194
rect 509 86 543 120
rect 609 176 643 210
rect 609 86 643 120
rect 695 176 729 210
rect 695 86 729 120
<< pdiffc >>
rect 83 522 117 556
rect 83 451 117 485
rect 83 380 117 414
rect 281 522 315 556
rect 281 451 315 485
rect 281 380 315 414
rect 409 548 443 582
rect 409 480 443 514
rect 409 412 443 446
rect 509 546 543 580
rect 509 463 543 497
rect 509 380 543 414
rect 609 546 643 580
rect 609 428 643 462
<< poly >>
rect 127 568 163 594
rect 211 568 247 594
rect 325 568 361 594
rect 463 592 499 618
rect 553 592 589 618
rect 127 310 163 368
rect 21 294 163 310
rect 21 260 37 294
rect 71 260 105 294
rect 139 280 163 294
rect 211 310 247 368
rect 325 310 361 368
rect 463 310 499 368
rect 553 322 589 368
rect 553 310 593 322
rect 211 294 277 310
rect 139 260 155 280
rect 21 244 155 260
rect 211 260 227 294
rect 261 260 277 294
rect 211 244 277 260
rect 325 294 391 310
rect 325 260 341 294
rect 375 260 391 294
rect 325 244 391 260
rect 463 294 593 310
rect 463 260 479 294
rect 513 274 593 294
rect 513 260 684 274
rect 463 244 684 260
rect 125 222 155 244
rect 247 222 277 244
rect 342 222 372 244
rect 568 222 598 244
rect 654 222 684 244
rect 125 48 155 74
rect 247 48 277 74
rect 342 48 372 74
rect 568 48 598 74
rect 654 48 684 74
<< polycont >>
rect 37 260 71 294
rect 105 260 139 294
rect 227 260 261 294
rect 341 260 375 294
rect 479 260 513 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 67 556 133 649
rect 393 582 459 649
rect 67 522 83 556
rect 117 522 133 556
rect 67 485 133 522
rect 67 451 83 485
rect 117 451 133 485
rect 67 414 133 451
rect 67 380 83 414
rect 117 380 133 414
rect 67 364 133 380
rect 265 556 331 572
rect 265 522 281 556
rect 315 522 331 556
rect 265 485 331 522
rect 265 451 281 485
rect 315 451 331 485
rect 265 414 331 451
rect 265 380 281 414
rect 315 380 331 414
rect 393 548 409 582
rect 443 548 459 582
rect 393 514 459 548
rect 393 480 409 514
rect 443 480 459 514
rect 393 446 459 480
rect 393 412 409 446
rect 443 412 459 446
rect 493 580 559 596
rect 493 546 509 580
rect 543 546 559 580
rect 493 497 559 546
rect 493 463 509 497
rect 543 463 559 497
rect 493 414 559 463
rect 265 378 331 380
rect 493 380 509 414
rect 543 380 559 414
rect 593 580 659 649
rect 593 546 609 580
rect 643 546 659 580
rect 593 462 659 546
rect 593 428 609 462
rect 643 428 659 462
rect 593 412 659 428
rect 493 378 559 380
rect 265 344 459 378
rect 493 344 659 378
rect 425 310 459 344
rect 21 294 167 310
rect 21 260 37 294
rect 71 260 105 294
rect 139 260 167 294
rect 21 236 167 260
rect 211 294 277 310
rect 211 260 227 294
rect 261 260 277 294
rect 211 236 277 260
rect 313 294 391 310
rect 313 260 341 294
rect 375 260 391 294
rect 313 236 391 260
rect 425 294 529 310
rect 425 260 479 294
rect 513 260 529 294
rect 425 244 529 260
rect 425 202 459 244
rect 593 210 659 344
rect 50 168 66 202
rect 100 168 297 202
rect 331 168 347 202
rect 50 118 116 168
rect 50 84 66 118
rect 100 84 116 118
rect 50 68 116 84
rect 150 86 181 120
rect 215 86 247 120
rect 150 17 247 86
rect 281 118 347 168
rect 281 84 297 118
rect 331 84 347 118
rect 281 68 347 84
rect 381 186 459 202
rect 381 152 383 186
rect 417 152 459 186
rect 381 118 459 152
rect 381 84 383 118
rect 417 84 459 118
rect 381 68 459 84
rect 493 194 559 210
rect 493 160 509 194
rect 543 160 559 194
rect 493 120 559 160
rect 493 86 509 120
rect 543 86 559 120
rect 493 17 559 86
rect 593 176 609 210
rect 643 176 659 210
rect 593 120 659 176
rect 593 86 609 120
rect 643 86 659 120
rect 593 70 659 86
rect 695 210 745 226
rect 729 176 745 210
rect 695 120 745 176
rect 729 86 745 120
rect 695 17 745 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 o21a_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 1034154
string GDS_START 1027326
<< end >>
