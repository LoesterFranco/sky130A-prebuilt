magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 95 196 161 398
rect 263 236 355 310
rect 2231 430 2293 596
rect 2137 364 2293 430
rect 2259 226 2293 364
rect 2220 70 2293 226
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 23 472 73 596
rect 113 506 179 649
rect 315 506 381 649
rect 421 578 759 612
rect 421 480 455 578
rect 23 446 359 472
rect 489 452 589 544
rect 623 452 691 544
rect 489 446 523 452
rect 23 438 523 446
rect 23 153 57 438
rect 325 412 523 438
rect 195 378 291 404
rect 195 344 455 378
rect 195 202 229 344
rect 389 260 455 344
rect 23 79 73 153
rect 109 17 159 153
rect 195 70 287 202
rect 323 17 373 202
rect 409 85 443 226
rect 489 185 523 412
rect 557 276 623 410
rect 489 119 555 185
rect 589 85 623 276
rect 409 51 623 85
rect 657 242 691 452
rect 725 482 759 578
rect 814 582 848 649
rect 814 516 915 582
rect 949 578 1138 612
rect 949 482 983 578
rect 725 448 983 482
rect 1017 464 1070 544
rect 1104 498 1138 578
rect 1172 532 1222 649
rect 1364 546 1494 596
rect 1364 510 1586 546
rect 1620 544 1686 649
rect 1726 510 1776 596
rect 1822 532 1888 649
rect 1104 464 1317 498
rect 725 276 783 448
rect 1017 414 1051 464
rect 846 348 1051 414
rect 1085 424 1223 430
rect 1085 390 1183 424
rect 1217 390 1223 424
rect 1085 358 1223 390
rect 817 280 1249 314
rect 817 242 851 280
rect 657 208 851 242
rect 885 210 954 246
rect 990 244 1249 280
rect 1183 243 1249 244
rect 1283 290 1317 464
rect 1364 358 1414 510
rect 1552 498 1776 510
rect 1458 430 1518 476
rect 1552 464 1894 498
rect 1458 396 1532 430
rect 1364 324 1464 358
rect 1283 224 1392 290
rect 657 80 723 208
rect 885 176 1032 210
rect 854 17 920 142
rect 954 114 1032 176
rect 1130 17 1249 206
rect 1283 90 1317 224
rect 1430 190 1464 324
rect 1365 124 1464 190
rect 1498 90 1532 396
rect 1566 248 1629 426
rect 1663 424 1746 430
rect 1697 390 1746 424
rect 1663 296 1746 390
rect 1828 323 1894 464
rect 1928 248 1978 596
rect 1566 214 1978 248
rect 1283 56 1532 90
rect 1705 17 1872 180
rect 1906 127 1978 214
rect 2018 326 2090 572
rect 2131 464 2197 649
rect 2327 364 2377 649
rect 2018 260 2225 326
rect 2018 90 2084 260
rect 2120 17 2186 226
rect 2327 17 2377 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 1183 390 1217 424
rect 1663 390 1697 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 1171 424 1229 430
rect 1171 390 1183 424
rect 1217 421 1229 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 1217 393 1663 421
rect 1217 390 1229 393
rect 1171 384 1229 390
rect 1651 390 1663 393
rect 1697 390 1709 424
rect 1651 384 1709 390
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
rlabel locali s 95 196 161 398 6 D
port 1 nsew signal input
rlabel locali s 2259 226 2293 364 6 Q
port 2 nsew signal output
rlabel locali s 2231 430 2293 596 6 Q
port 2 nsew signal output
rlabel locali s 2220 70 2293 226 6 Q
port 2 nsew signal output
rlabel locali s 2137 364 2293 430 6 Q
port 2 nsew signal output
rlabel metal1 s 1651 421 1709 430 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1651 384 1709 393 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1171 421 1229 430 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1171 393 1709 421 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1171 384 1229 393 6 SET_B
port 3 nsew signal input
rlabel locali s 263 236 355 310 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2400 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 2400 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2732390
string GDS_START 2715206
<< end >>
