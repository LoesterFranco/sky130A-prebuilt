magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1196 561
rect 457 455 523 527
rect 629 455 695 527
rect 801 455 867 527
rect 973 455 1039 527
rect 116 341 349 407
rect 116 317 376 341
rect 18 207 286 283
rect 18 199 80 207
rect 320 179 376 317
rect 410 296 1094 341
rect 410 213 479 296
rect 513 213 800 262
rect 845 215 1094 296
rect 320 173 781 179
rect 18 17 85 161
rect 119 139 781 173
rect 119 123 329 139
rect 455 135 781 139
rect 119 74 157 123
rect 191 17 257 89
rect 291 51 329 123
rect 367 17 423 105
rect 901 17 939 113
rect 1073 17 1125 177
rect 0 -17 1196 17
<< obsli1 >>
rect 36 443 423 493
rect 36 359 75 443
rect 191 441 423 443
rect 383 421 423 441
rect 557 421 595 493
rect 729 421 767 493
rect 901 421 937 493
rect 1073 421 1125 493
rect 383 375 1125 421
rect 815 147 1039 181
rect 815 101 867 147
rect 457 51 867 101
rect 973 51 1039 147
<< metal1 >>
rect 0 496 1196 592
rect 0 -48 1196 48
<< labels >>
rlabel locali s 513 213 800 262 6 A1
port 1 nsew signal input
rlabel locali s 845 215 1094 296 6 A2
port 2 nsew signal input
rlabel locali s 410 296 1094 341 6 A2
port 2 nsew signal input
rlabel locali s 410 213 479 296 6 A2
port 2 nsew signal input
rlabel locali s 18 207 286 283 6 B1
port 3 nsew signal input
rlabel locali s 18 199 80 207 6 B1
port 3 nsew signal input
rlabel locali s 455 135 781 139 6 Y
port 4 nsew signal output
rlabel locali s 320 179 376 317 6 Y
port 4 nsew signal output
rlabel locali s 320 173 781 179 6 Y
port 4 nsew signal output
rlabel locali s 291 51 329 123 6 Y
port 4 nsew signal output
rlabel locali s 119 139 781 173 6 Y
port 4 nsew signal output
rlabel locali s 119 123 329 139 6 Y
port 4 nsew signal output
rlabel locali s 119 74 157 123 6 Y
port 4 nsew signal output
rlabel locali s 116 341 349 407 6 Y
port 4 nsew signal output
rlabel locali s 116 317 376 341 6 Y
port 4 nsew signal output
rlabel locali s 1073 17 1125 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 901 17 939 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 367 17 423 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 191 17 257 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 18 17 85 161 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1196 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 973 455 1039 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 801 455 867 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 629 455 695 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 457 455 523 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1196 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4058102
string GDS_START 4049568
<< end >>
