magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 123 424 273 596
rect 407 424 473 596
rect 792 424 858 596
rect 25 390 858 424
rect 25 236 71 390
rect 407 364 473 390
rect 792 364 858 390
rect 105 270 307 356
rect 512 326 743 356
rect 899 326 1223 356
rect 426 270 743 326
rect 828 268 1223 326
rect 25 202 345 236
rect 107 119 173 202
rect 279 119 345 202
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 458 89 649
rect 307 458 373 649
rect 507 458 758 649
rect 892 390 1153 649
rect 21 85 71 168
rect 209 85 243 168
rect 381 85 415 234
rect 451 184 1125 234
rect 451 119 517 184
rect 551 85 589 150
rect 623 119 689 184
rect 723 85 775 150
rect 21 51 775 85
rect 817 17 883 150
rect 917 78 955 184
rect 989 17 1055 150
rect 1091 78 1125 184
rect 1161 17 1227 234
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 105 270 307 356 6 A
port 1 nsew signal input
rlabel locali s 512 326 743 356 6 B
port 2 nsew signal input
rlabel locali s 426 270 743 326 6 B
port 2 nsew signal input
rlabel locali s 899 326 1223 356 6 C
port 3 nsew signal input
rlabel locali s 828 268 1223 326 6 C
port 3 nsew signal input
rlabel locali s 792 424 858 596 6 Y
port 4 nsew signal output
rlabel locali s 792 364 858 390 6 Y
port 4 nsew signal output
rlabel locali s 407 424 473 596 6 Y
port 4 nsew signal output
rlabel locali s 407 364 473 390 6 Y
port 4 nsew signal output
rlabel locali s 279 119 345 202 6 Y
port 4 nsew signal output
rlabel locali s 123 424 273 596 6 Y
port 4 nsew signal output
rlabel locali s 107 119 173 202 6 Y
port 4 nsew signal output
rlabel locali s 25 390 858 424 6 Y
port 4 nsew signal output
rlabel locali s 25 236 71 390 6 Y
port 4 nsew signal output
rlabel locali s 25 202 345 236 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1248 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2099546
string GDS_START 2088846
<< end >>
