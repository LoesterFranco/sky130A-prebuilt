magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 644 561
rect 110 435 153 527
rect 17 211 111 323
rect 382 383 454 527
rect 488 299 540 493
rect 110 17 153 109
rect 506 165 540 299
rect 382 17 448 113
rect 482 51 540 165
rect 0 -17 644 17
<< obsli1 >>
rect 17 401 76 493
rect 187 435 264 493
rect 17 357 179 401
rect 145 265 179 357
rect 145 199 196 265
rect 230 255 264 435
rect 303 349 348 486
rect 303 315 448 349
rect 414 265 448 315
rect 230 215 380 255
rect 145 177 179 199
rect 19 143 179 177
rect 19 51 76 143
rect 230 109 264 215
rect 414 199 472 265
rect 414 181 448 199
rect 187 51 264 109
rect 303 147 448 181
rect 303 51 348 147
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 17 211 111 323 6 A
port 1 nsew signal input
rlabel locali s 506 165 540 299 6 X
port 2 nsew signal output
rlabel locali s 488 299 540 493 6 X
port 2 nsew signal output
rlabel locali s 482 51 540 165 6 X
port 2 nsew signal output
rlabel locali s 382 17 448 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 110 17 153 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 644 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 382 383 454 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 110 435 153 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 644 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 644 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2811608
string GDS_START 2806206
<< end >>
