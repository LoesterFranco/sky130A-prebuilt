magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 552 561
rect 19 299 85 527
rect 17 149 85 265
rect 119 259 191 493
rect 231 293 297 527
rect 337 259 403 493
rect 443 293 509 527
rect 119 203 403 259
rect 119 136 191 203
rect 19 17 85 115
rect 119 51 243 136
rect 335 17 401 155
rect 0 -17 552 17
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 17 149 85 265 6 A
port 1 nsew signal input
rlabel locali s 337 259 403 493 6 Y
port 2 nsew signal output
rlabel locali s 119 259 191 493 6 Y
port 2 nsew signal output
rlabel locali s 119 203 403 259 6 Y
port 2 nsew signal output
rlabel locali s 119 136 191 203 6 Y
port 2 nsew signal output
rlabel locali s 119 51 243 136 6 Y
port 2 nsew signal output
rlabel locali s 335 17 401 155 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 19 17 85 115 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 443 293 509 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 231 293 297 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 19 299 85 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 552 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3243348
string GDS_START 3238308
<< end >>
