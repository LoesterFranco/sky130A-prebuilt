magic
tech sky130A
magscale 1 2
timestamp 1601050039
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 257 47 287 177
rect 341 47 371 177
<< pmoshvt >>
rect 89 297 119 497
rect 173 297 203 497
rect 257 297 287 497
rect 341 297 371 497
<< ndiff >>
rect 37 93 89 177
rect 37 59 45 93
rect 79 59 89 93
rect 37 47 89 59
rect 119 101 173 177
rect 119 67 129 101
rect 163 67 173 101
rect 119 47 173 67
rect 203 93 257 177
rect 203 59 213 93
rect 247 59 257 93
rect 203 47 257 59
rect 287 101 341 177
rect 287 67 297 101
rect 331 67 341 101
rect 287 47 341 67
rect 371 94 423 177
rect 371 60 381 94
rect 415 60 423 94
rect 371 47 423 60
<< pdiff >>
rect 37 485 89 497
rect 37 451 45 485
rect 79 451 89 485
rect 37 417 89 451
rect 37 383 45 417
rect 79 383 89 417
rect 37 349 89 383
rect 37 315 45 349
rect 79 315 89 349
rect 37 297 89 315
rect 119 485 173 497
rect 119 451 129 485
rect 163 451 173 485
rect 119 417 173 451
rect 119 383 129 417
rect 163 383 173 417
rect 119 349 173 383
rect 119 315 129 349
rect 163 315 173 349
rect 119 297 173 315
rect 203 485 257 497
rect 203 451 213 485
rect 247 451 257 485
rect 203 417 257 451
rect 203 383 213 417
rect 247 383 257 417
rect 203 297 257 383
rect 287 485 341 497
rect 287 451 297 485
rect 331 451 341 485
rect 287 417 341 451
rect 287 383 297 417
rect 331 383 341 417
rect 287 349 341 383
rect 287 315 297 349
rect 331 315 341 349
rect 287 297 341 315
rect 371 485 423 497
rect 371 451 381 485
rect 415 451 423 485
rect 371 297 423 451
<< ndiffc >>
rect 45 59 79 93
rect 129 67 163 101
rect 213 59 247 93
rect 297 67 331 101
rect 381 60 415 94
<< pdiffc >>
rect 45 451 79 485
rect 45 383 79 417
rect 45 315 79 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 213 451 247 485
rect 213 383 247 417
rect 297 451 331 485
rect 297 383 331 417
rect 297 315 331 349
rect 381 451 415 485
<< poly >>
rect 89 497 119 523
rect 173 497 203 523
rect 257 497 287 523
rect 341 497 371 523
rect 89 265 119 297
rect 173 265 203 297
rect 257 265 287 297
rect 341 265 371 297
rect 21 249 371 265
rect 21 215 37 249
rect 71 215 129 249
rect 163 215 213 249
rect 247 215 297 249
rect 331 215 371 249
rect 21 199 371 215
rect 89 177 119 199
rect 173 177 203 199
rect 257 177 287 199
rect 341 177 371 199
rect 89 21 119 47
rect 173 21 203 47
rect 257 21 287 47
rect 341 21 371 47
<< polycont >>
rect 37 215 71 249
rect 129 215 163 249
rect 213 215 247 249
rect 297 215 331 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 26 485 79 527
rect 26 451 45 485
rect 26 417 79 451
rect 26 383 45 417
rect 26 349 79 383
rect 26 315 45 349
rect 26 299 79 315
rect 113 485 179 493
rect 113 451 129 485
rect 163 451 179 485
rect 113 417 179 451
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 213 485 247 527
rect 213 417 247 451
rect 213 367 247 383
rect 281 485 347 493
rect 281 451 297 485
rect 331 451 347 485
rect 281 417 347 451
rect 381 485 423 527
rect 415 451 423 485
rect 381 435 423 451
rect 281 383 297 417
rect 331 383 347 417
rect 113 315 129 349
rect 163 333 179 349
rect 281 349 347 383
rect 281 333 297 349
rect 163 315 297 333
rect 331 337 347 349
rect 331 315 434 337
rect 113 299 434 315
rect 21 249 347 265
rect 21 215 37 249
rect 71 215 129 249
rect 163 215 213 249
rect 247 215 297 249
rect 331 215 347 249
rect 381 181 434 299
rect 113 145 434 181
rect 26 93 79 109
rect 26 59 45 93
rect 26 17 79 59
rect 113 101 179 145
rect 113 67 129 101
rect 163 67 179 101
rect 113 51 179 67
rect 213 93 247 109
rect 213 17 247 59
rect 281 101 347 145
rect 281 67 297 101
rect 331 67 347 101
rect 281 51 347 67
rect 381 94 431 110
rect 415 60 431 94
rect 381 17 431 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel corelocali s 397 153 431 187 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 397 289 431 323 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 121 221 155 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 213 221 247 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 305 221 339 255 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
rlabel comment s 0 0 0 0 4 inv_4
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2235240
string GDS_START 2230250
string path 0.000 0.000 11.500 0.000 
<< end >>
