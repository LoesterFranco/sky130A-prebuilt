magic
tech sky130A
magscale 1 2
timestamp 1601050058
<< locali >>
rect 703 393 753 425
rect 871 393 921 425
rect 703 391 921 393
rect 1123 391 1179 493
rect 703 357 1179 391
rect 703 289 1033 323
rect 703 257 737 289
rect 18 215 365 257
rect 419 215 737 257
rect 999 257 1033 289
rect 771 215 953 255
rect 999 215 1083 257
rect 1121 181 1179 357
rect 107 145 1179 181
rect 107 51 173 145
rect 275 51 341 145
rect 443 51 509 145
rect 611 51 677 145
rect 779 51 845 145
rect 947 51 1013 145
rect 1121 51 1179 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 30 325 81 493
rect 115 359 165 527
rect 199 325 249 493
rect 283 359 333 527
rect 367 417 585 493
rect 367 325 417 417
rect 30 291 417 325
rect 451 325 501 383
rect 535 359 585 417
rect 619 459 1005 493
rect 619 325 669 459
rect 787 427 837 459
rect 955 427 1005 459
rect 1039 425 1089 493
rect 451 291 669 325
rect 18 17 73 181
rect 207 17 241 111
rect 375 17 409 111
rect 543 17 577 111
rect 711 17 745 111
rect 879 17 913 111
rect 1047 17 1081 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< obsm1 >>
rect 477 456 536 467
rect 1029 456 1088 467
rect 477 428 1088 456
rect 477 413 536 428
rect 1029 413 1088 428
<< labels >>
rlabel locali s 18 215 365 257 6 A
port 1 nsew signal input
rlabel locali s 999 257 1033 289 6 B
port 2 nsew signal input
rlabel locali s 999 215 1083 257 6 B
port 2 nsew signal input
rlabel locali s 703 289 1033 323 6 B
port 2 nsew signal input
rlabel locali s 703 257 737 289 6 B
port 2 nsew signal input
rlabel locali s 419 215 737 257 6 B
port 2 nsew signal input
rlabel locali s 771 215 953 255 6 C
port 3 nsew signal input
rlabel locali s 1123 391 1179 493 6 Y
port 4 nsew signal output
rlabel locali s 1121 181 1179 357 6 Y
port 4 nsew signal output
rlabel locali s 1121 51 1179 145 6 Y
port 4 nsew signal output
rlabel locali s 947 51 1013 145 6 Y
port 4 nsew signal output
rlabel locali s 871 393 921 425 6 Y
port 4 nsew signal output
rlabel locali s 779 51 845 145 6 Y
port 4 nsew signal output
rlabel locali s 703 393 753 425 6 Y
port 4 nsew signal output
rlabel locali s 703 391 921 393 6 Y
port 4 nsew signal output
rlabel locali s 703 357 1179 391 6 Y
port 4 nsew signal output
rlabel locali s 611 51 677 145 6 Y
port 4 nsew signal output
rlabel locali s 443 51 509 145 6 Y
port 4 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 4 nsew signal output
rlabel locali s 107 145 1179 181 6 Y
port 4 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1988588
string GDS_START 1979272
<< end >>
