magic
tech sky130A
magscale 1 2
timestamp 1601050056
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 227 368 263 536
rect 317 368 353 536
rect 407 368 443 536
rect 524 368 560 592
<< nmoslvt >>
rect 84 74 114 184
rect 323 98 353 226
rect 401 98 431 226
rect 558 78 588 226
<< ndiff >>
rect 266 214 323 226
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 136 185 184
rect 114 102 139 136
rect 173 102 185 136
rect 114 74 185 102
rect 266 180 278 214
rect 312 180 323 214
rect 266 144 323 180
rect 266 110 278 144
rect 312 110 323 144
rect 266 98 323 110
rect 353 98 401 226
rect 431 146 558 226
rect 431 112 442 146
rect 476 112 513 146
rect 547 112 558 146
rect 431 98 558 112
rect 508 78 558 98
rect 588 214 645 226
rect 588 180 599 214
rect 633 180 645 214
rect 588 124 645 180
rect 588 90 599 124
rect 633 90 645 124
rect 588 78 645 90
<< pdiff >>
rect 458 576 524 592
rect 458 542 470 576
rect 504 542 524 576
rect 458 536 524 542
rect 27 514 227 536
rect 27 480 39 514
rect 73 480 111 514
rect 145 480 183 514
rect 217 480 227 514
rect 27 368 227 480
rect 263 524 317 536
rect 263 490 273 524
rect 307 490 317 524
rect 263 414 317 490
rect 263 380 273 414
rect 307 380 317 414
rect 263 368 317 380
rect 353 524 407 536
rect 353 490 363 524
rect 397 490 407 524
rect 353 440 407 490
rect 353 406 363 440
rect 397 406 407 440
rect 353 368 407 406
rect 443 504 524 536
rect 443 470 470 504
rect 504 470 524 504
rect 443 426 524 470
rect 443 392 470 426
rect 504 392 524 426
rect 443 368 524 392
rect 560 580 616 592
rect 560 546 570 580
rect 604 546 616 580
rect 560 497 616 546
rect 560 463 570 497
rect 604 463 616 497
rect 560 414 616 463
rect 560 380 570 414
rect 604 380 616 414
rect 560 368 616 380
<< ndiffc >>
rect 39 112 73 146
rect 139 102 173 136
rect 278 180 312 214
rect 278 110 312 144
rect 442 112 476 146
rect 513 112 547 146
rect 599 180 633 214
rect 599 90 633 124
<< pdiffc >>
rect 470 542 504 576
rect 39 480 73 514
rect 111 480 145 514
rect 183 480 217 514
rect 273 490 307 524
rect 273 380 307 414
rect 363 490 397 524
rect 363 406 397 440
rect 470 470 504 504
rect 470 392 504 426
rect 570 546 604 580
rect 570 463 604 497
rect 570 380 604 414
<< poly >>
rect 524 592 560 618
rect 227 536 263 562
rect 317 536 353 562
rect 407 536 443 562
rect 227 350 263 368
rect 44 320 263 350
rect 44 286 60 320
rect 94 286 114 320
rect 44 270 114 286
rect 317 272 353 368
rect 407 336 443 368
rect 84 184 114 270
rect 162 256 353 272
rect 162 222 178 256
rect 212 242 353 256
rect 212 222 228 242
rect 323 226 353 242
rect 401 320 475 336
rect 524 330 560 368
rect 401 286 425 320
rect 459 286 475 320
rect 401 270 475 286
rect 517 314 588 330
rect 517 280 533 314
rect 567 280 588 314
rect 401 226 431 270
rect 517 264 588 280
rect 558 226 588 264
rect 162 206 228 222
rect 84 48 114 74
rect 323 72 353 98
rect 401 72 431 98
rect 558 52 588 78
<< polycont >>
rect 60 286 94 320
rect 178 222 212 256
rect 425 286 459 320
rect 533 280 567 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 514 233 530
rect 23 480 39 514
rect 73 480 111 514
rect 145 480 183 514
rect 217 480 233 514
rect 23 464 233 480
rect 273 524 307 649
rect 454 576 520 649
rect 454 542 470 576
rect 504 542 520 576
rect 25 320 110 430
rect 25 286 60 320
rect 94 286 110 320
rect 25 270 110 286
rect 162 256 228 464
rect 273 414 307 490
rect 273 364 307 380
rect 341 524 413 540
rect 341 490 363 524
rect 397 490 413 524
rect 341 440 413 490
rect 341 406 363 440
rect 397 406 413 440
rect 341 390 413 406
rect 454 504 520 542
rect 454 470 470 504
rect 504 470 520 504
rect 454 426 520 470
rect 454 392 470 426
rect 504 392 520 426
rect 454 390 520 392
rect 554 580 651 596
rect 554 546 570 580
rect 604 546 651 580
rect 554 497 651 546
rect 554 463 570 497
rect 604 463 651 497
rect 554 414 651 463
rect 162 236 178 256
rect 23 222 178 236
rect 212 222 228 256
rect 341 230 375 390
rect 554 380 570 414
rect 604 380 651 414
rect 554 364 651 380
rect 409 320 475 356
rect 409 286 425 320
rect 459 286 475 320
rect 409 270 475 286
rect 515 314 583 330
rect 515 280 533 314
rect 567 280 583 314
rect 515 264 583 280
rect 515 230 549 264
rect 617 230 651 364
rect 23 202 228 222
rect 262 214 549 230
rect 23 146 89 202
rect 262 180 278 214
rect 312 196 549 214
rect 583 214 651 230
rect 312 180 328 196
rect 23 112 39 146
rect 73 112 89 146
rect 23 70 89 112
rect 123 136 189 168
rect 123 102 139 136
rect 173 102 189 136
rect 123 17 189 102
rect 262 144 328 180
rect 583 180 599 214
rect 633 180 651 214
rect 262 110 278 144
rect 312 110 328 144
rect 262 94 328 110
rect 426 146 549 162
rect 426 112 442 146
rect 476 112 513 146
rect 547 112 549 146
rect 426 17 549 112
rect 583 124 651 180
rect 583 90 599 124
rect 633 90 651 124
rect 583 74 651 90
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 and2b_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 7 nsew
flabel corelocali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 3196124
string GDS_START 3190134
<< end >>
