magic
tech sky130A
magscale 1 2
timestamp 1601050088
<< locali >>
rect 537 390 1170 428
rect 85 270 219 356
rect 750 364 1170 390
rect 353 270 647 356
rect 985 226 1031 364
rect 1164 236 1415 330
rect 826 160 1069 226
rect 985 154 1069 160
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 458 89 649
rect 298 530 513 649
rect 627 530 726 649
rect 916 530 1080 649
rect 1194 530 1513 649
rect 123 462 1246 496
rect 123 424 157 462
rect 17 390 157 424
rect 191 390 287 428
rect 17 150 51 390
rect 253 236 287 390
rect 1212 398 1246 462
rect 1280 432 1513 530
rect 1212 364 1483 398
rect 720 260 922 326
rect 720 236 754 260
rect 85 202 754 236
rect 85 184 151 202
rect 292 150 594 168
rect 17 134 594 150
rect 17 116 358 134
rect 187 17 256 82
rect 292 78 358 116
rect 394 17 492 100
rect 528 78 594 134
rect 628 17 694 168
rect 1449 202 1483 364
rect 1189 168 1483 202
rect 740 120 806 126
rect 1103 120 1513 134
rect 740 70 1513 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
rlabel locali s 85 270 219 356 6 A_N
port 1 nsew signal input
rlabel locali s 1164 236 1415 330 6 B
port 2 nsew signal input
rlabel locali s 353 270 647 356 6 C
port 3 nsew signal input
rlabel locali s 985 226 1031 364 6 Y
port 4 nsew signal output
rlabel locali s 985 154 1069 160 6 Y
port 4 nsew signal output
rlabel locali s 826 160 1069 226 6 Y
port 4 nsew signal output
rlabel locali s 750 364 1170 390 6 Y
port 4 nsew signal output
rlabel locali s 537 390 1170 428 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -49 1536 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 617 1536 715 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2066032
string GDS_START 2055924
<< end >>
