magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 583 323 659 493
rect 771 323 847 493
rect 959 323 1035 493
rect 1147 323 1223 493
rect 583 289 1361 323
rect 17 215 101 255
rect 1283 181 1361 289
rect 583 147 1361 181
rect 583 52 659 147
rect 771 52 847 147
rect 959 52 1035 147
rect 1147 52 1223 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 289 69 527
rect 103 309 179 493
rect 145 255 179 309
rect 217 323 283 493
rect 327 357 361 527
rect 395 323 471 493
rect 515 357 549 527
rect 703 367 737 527
rect 891 367 925 527
rect 1079 367 1113 527
rect 1267 367 1301 527
rect 217 289 549 323
rect 515 255 549 289
rect 145 215 471 255
rect 515 215 1249 255
rect 145 181 179 215
rect 515 181 549 215
rect 35 17 69 181
rect 103 52 179 181
rect 217 147 549 181
rect 217 52 283 147
rect 327 17 361 113
rect 395 52 471 147
rect 515 17 549 113
rect 703 17 737 113
rect 891 17 925 113
rect 1079 17 1113 113
rect 1267 17 1301 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
rlabel locali s 17 215 101 255 6 A
port 1 nsew signal input
rlabel locali s 1283 181 1361 289 6 Y
port 2 nsew signal output
rlabel locali s 1147 323 1223 493 6 Y
port 2 nsew signal output
rlabel locali s 1147 52 1223 147 6 Y
port 2 nsew signal output
rlabel locali s 959 323 1035 493 6 Y
port 2 nsew signal output
rlabel locali s 959 52 1035 147 6 Y
port 2 nsew signal output
rlabel locali s 771 323 847 493 6 Y
port 2 nsew signal output
rlabel locali s 771 52 847 147 6 Y
port 2 nsew signal output
rlabel locali s 583 323 659 493 6 Y
port 2 nsew signal output
rlabel locali s 583 289 1361 323 6 Y
port 2 nsew signal output
rlabel locali s 583 147 1361 181 6 Y
port 2 nsew signal output
rlabel locali s 583 52 659 147 6 Y
port 2 nsew signal output
rlabel metal1 s 0 -48 1380 48 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1743172
string GDS_START 1732476
<< end >>
