magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 81 74 111 222
rect 167 74 197 222
rect 361 74 391 222
rect 461 74 491 222
rect 541 74 571 222
rect 649 74 679 222
<< pmoshvt >>
rect 160 368 190 592
rect 250 368 280 592
rect 358 368 388 568
rect 448 368 478 568
rect 548 368 578 568
rect 652 368 682 568
<< ndiff >>
rect 28 210 81 222
rect 28 176 36 210
rect 70 176 81 210
rect 28 120 81 176
rect 28 86 36 120
rect 70 86 81 120
rect 28 74 81 86
rect 111 210 167 222
rect 111 176 122 210
rect 156 176 167 210
rect 111 120 167 176
rect 111 86 122 120
rect 156 86 167 120
rect 111 74 167 86
rect 197 152 250 222
rect 197 118 208 152
rect 242 118 250 152
rect 197 74 250 118
rect 304 152 361 222
rect 304 118 316 152
rect 350 118 361 152
rect 304 74 361 118
rect 391 169 461 222
rect 391 135 416 169
rect 450 135 461 169
rect 391 74 461 135
rect 491 74 541 222
rect 571 152 649 222
rect 571 118 590 152
rect 624 118 649 152
rect 571 74 649 118
rect 679 210 736 222
rect 679 176 690 210
rect 724 176 736 210
rect 679 120 736 176
rect 679 86 690 120
rect 724 86 736 120
rect 679 74 736 86
<< pdiff >>
rect 105 580 160 592
rect 105 546 113 580
rect 147 546 160 580
rect 105 462 160 546
rect 105 428 113 462
rect 147 428 160 462
rect 105 368 160 428
rect 190 580 250 592
rect 190 546 203 580
rect 237 546 250 580
rect 190 508 250 546
rect 190 474 203 508
rect 237 474 250 508
rect 190 368 250 474
rect 280 568 333 592
rect 280 560 358 568
rect 280 526 293 560
rect 327 526 358 560
rect 280 492 358 526
rect 280 458 293 492
rect 327 458 358 492
rect 280 368 358 458
rect 388 560 448 568
rect 388 526 401 560
rect 435 526 448 560
rect 388 492 448 526
rect 388 458 401 492
rect 435 458 448 492
rect 388 368 448 458
rect 478 531 548 568
rect 478 497 491 531
rect 525 497 548 531
rect 478 440 548 497
rect 478 406 491 440
rect 525 406 548 440
rect 478 368 548 406
rect 578 560 652 568
rect 578 526 593 560
rect 627 526 652 560
rect 578 492 652 526
rect 578 458 593 492
rect 627 458 652 492
rect 578 424 652 458
rect 578 390 593 424
rect 627 390 652 424
rect 578 368 652 390
rect 682 556 737 568
rect 682 522 695 556
rect 729 522 737 556
rect 682 440 737 522
rect 682 406 695 440
rect 729 406 737 440
rect 682 368 737 406
<< ndiffc >>
rect 36 176 70 210
rect 36 86 70 120
rect 122 176 156 210
rect 122 86 156 120
rect 208 118 242 152
rect 316 118 350 152
rect 416 135 450 169
rect 590 118 624 152
rect 690 176 724 210
rect 690 86 724 120
<< pdiffc >>
rect 113 546 147 580
rect 113 428 147 462
rect 203 546 237 580
rect 203 474 237 508
rect 293 526 327 560
rect 293 458 327 492
rect 401 526 435 560
rect 401 458 435 492
rect 491 497 525 531
rect 491 406 525 440
rect 593 526 627 560
rect 593 458 627 492
rect 593 390 627 424
rect 695 522 729 556
rect 695 406 729 440
<< poly >>
rect 160 592 190 618
rect 250 592 280 618
rect 358 568 388 594
rect 448 568 478 594
rect 548 568 578 594
rect 652 568 682 594
rect 160 353 190 368
rect 250 353 280 368
rect 358 353 388 368
rect 448 353 478 368
rect 548 353 578 368
rect 652 353 682 368
rect 157 310 193 353
rect 247 310 283 353
rect 355 336 391 353
rect 445 336 481 353
rect 545 336 581 353
rect 649 336 685 353
rect 81 294 283 310
rect 81 260 233 294
rect 267 260 283 294
rect 325 320 391 336
rect 325 286 341 320
rect 375 286 391 320
rect 325 270 391 286
rect 433 320 499 336
rect 433 286 449 320
rect 483 286 499 320
rect 433 270 499 286
rect 541 320 607 336
rect 541 286 557 320
rect 591 286 607 320
rect 541 270 607 286
rect 649 320 747 336
rect 649 286 697 320
rect 731 286 747 320
rect 649 270 747 286
rect 81 244 283 260
rect 81 222 111 244
rect 167 222 197 244
rect 361 222 391 270
rect 461 222 491 270
rect 541 222 571 270
rect 649 222 679 270
rect 81 48 111 74
rect 167 48 197 74
rect 361 48 391 74
rect 461 48 491 74
rect 541 48 571 74
rect 649 48 679 74
<< polycont >>
rect 233 260 267 294
rect 341 286 375 320
rect 449 286 483 320
rect 557 286 591 320
rect 697 286 731 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 97 580 147 649
rect 97 546 113 580
rect 97 462 147 546
rect 97 428 113 462
rect 97 412 147 428
rect 181 580 237 596
rect 181 546 203 580
rect 181 508 237 546
rect 181 474 203 508
rect 181 458 237 474
rect 277 560 343 649
rect 277 526 293 560
rect 327 526 343 560
rect 277 492 343 526
rect 277 458 293 492
rect 327 458 343 492
rect 385 581 645 615
rect 385 560 451 581
rect 385 526 401 560
rect 435 526 451 560
rect 575 560 645 581
rect 385 492 451 526
rect 385 458 401 492
rect 435 458 451 492
rect 491 531 541 547
rect 525 497 541 531
rect 181 378 215 458
rect 491 440 541 497
rect 106 344 215 378
rect 249 406 491 424
rect 525 406 541 440
rect 249 390 541 406
rect 575 526 593 560
rect 627 526 645 560
rect 575 492 645 526
rect 575 458 593 492
rect 627 458 645 492
rect 575 424 645 458
rect 575 390 593 424
rect 627 390 645 424
rect 679 556 745 649
rect 679 522 695 556
rect 729 522 745 556
rect 679 440 745 522
rect 679 406 695 440
rect 729 406 745 440
rect 679 390 745 406
rect 20 210 70 226
rect 20 176 36 210
rect 20 120 70 176
rect 20 86 36 120
rect 20 17 70 86
rect 106 210 172 344
rect 249 310 283 390
rect 106 176 122 210
rect 156 176 172 210
rect 217 294 283 310
rect 217 260 233 294
rect 267 260 283 294
rect 317 320 381 356
rect 317 286 341 320
rect 375 286 381 320
rect 317 270 381 286
rect 415 320 499 356
rect 415 286 449 320
rect 483 286 499 320
rect 415 270 499 286
rect 541 320 647 356
rect 541 286 557 320
rect 591 286 647 320
rect 541 270 647 286
rect 681 320 747 356
rect 681 286 697 320
rect 731 286 747 320
rect 681 270 747 286
rect 217 236 283 260
rect 217 202 466 236
rect 106 120 172 176
rect 400 169 466 202
rect 106 86 122 120
rect 156 86 172 120
rect 106 70 172 86
rect 208 152 258 168
rect 242 118 258 152
rect 208 17 258 118
rect 300 152 366 168
rect 300 118 316 152
rect 350 118 366 152
rect 400 135 416 169
rect 450 135 466 169
rect 400 119 466 135
rect 500 210 740 236
rect 500 202 690 210
rect 300 85 366 118
rect 500 85 534 202
rect 674 176 690 202
rect 724 176 740 210
rect 300 51 534 85
rect 574 152 640 168
rect 574 118 590 152
rect 624 118 640 152
rect 574 17 640 118
rect 674 120 740 176
rect 674 86 690 120
rect 724 86 740 120
rect 674 70 740 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a22o_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3456310
string GDS_START 3449082
<< end >>
