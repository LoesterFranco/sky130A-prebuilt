magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 2726 704
rect 1629 311 1933 332
<< pwell >>
rect 0 0 2688 49
<< scpmos >>
rect 86 464 116 592
rect 186 464 216 592
rect 270 464 300 592
rect 508 464 538 592
rect 592 464 622 592
rect 706 464 736 592
rect 914 368 944 592
rect 1004 368 1034 592
rect 1212 457 1242 541
rect 1313 461 1343 545
rect 1397 461 1427 545
rect 1522 461 1552 545
rect 1724 347 1754 547
rect 1814 347 1844 547
rect 1963 508 1993 592
rect 2047 508 2077 592
rect 2162 508 2192 592
rect 2252 508 2282 592
rect 2369 424 2399 592
rect 2571 368 2601 592
<< nmoslvt >>
rect 84 88 114 172
rect 282 81 312 165
rect 360 81 390 165
rect 515 81 545 165
rect 593 81 623 165
rect 716 81 746 165
rect 918 74 948 222
rect 1005 74 1035 222
rect 1203 118 1233 202
rect 1289 118 1319 202
rect 1367 118 1397 202
rect 1445 118 1475 202
rect 1629 74 1659 202
rect 1715 74 1745 202
rect 1942 74 1972 158
rect 2014 74 2044 158
rect 2105 74 2135 158
rect 2177 74 2207 158
rect 2376 74 2406 184
rect 2574 74 2604 222
<< ndiff >>
rect 27 147 84 172
rect 27 113 39 147
rect 73 113 84 147
rect 27 88 84 113
rect 114 147 171 172
rect 861 202 918 222
rect 861 168 873 202
rect 907 168 918 202
rect 114 113 125 147
rect 159 113 171 147
rect 114 88 171 113
rect 225 127 282 165
rect 225 93 237 127
rect 271 93 282 127
rect 225 81 282 93
rect 312 81 360 165
rect 390 153 515 165
rect 390 119 470 153
rect 504 119 515 153
rect 390 81 515 119
rect 545 81 593 165
rect 623 127 716 165
rect 623 93 652 127
rect 686 93 716 127
rect 623 81 716 93
rect 746 130 803 165
rect 746 96 757 130
rect 791 96 803 130
rect 746 81 803 96
rect 861 120 918 168
rect 861 86 873 120
rect 907 86 918 120
rect 861 74 918 86
rect 948 127 1005 222
rect 948 93 959 127
rect 993 93 1005 127
rect 948 74 1005 93
rect 1035 210 1092 222
rect 1035 176 1046 210
rect 1080 176 1092 210
rect 1035 120 1092 176
rect 1035 86 1046 120
rect 1080 86 1092 120
rect 1146 179 1203 202
rect 1146 145 1158 179
rect 1192 145 1203 179
rect 1146 118 1203 145
rect 1233 179 1289 202
rect 1233 145 1244 179
rect 1278 145 1289 179
rect 1233 118 1289 145
rect 1319 118 1367 202
rect 1397 118 1445 202
rect 1475 118 1629 202
rect 1035 74 1092 86
rect 1490 82 1629 118
rect 1490 48 1502 82
rect 1536 74 1629 82
rect 1659 179 1715 202
rect 1659 145 1670 179
rect 1704 145 1715 179
rect 1659 74 1715 145
rect 1745 158 1795 202
rect 2517 210 2574 222
rect 1745 129 1942 158
rect 1745 95 1897 129
rect 1931 95 1942 129
rect 1745 74 1942 95
rect 1972 74 2014 158
rect 2044 133 2105 158
rect 2044 99 2055 133
rect 2089 99 2105 133
rect 2044 74 2105 99
rect 2135 74 2177 158
rect 2207 133 2264 158
rect 2207 99 2218 133
rect 2252 99 2264 133
rect 2207 74 2264 99
rect 2318 117 2376 184
rect 2318 83 2330 117
rect 2364 83 2376 117
rect 2318 74 2376 83
rect 2406 146 2463 184
rect 2406 112 2417 146
rect 2451 112 2463 146
rect 2406 74 2463 112
rect 2517 176 2529 210
rect 2563 176 2574 210
rect 2517 120 2574 176
rect 2517 86 2529 120
rect 2563 86 2574 120
rect 2517 74 2574 86
rect 2604 210 2661 222
rect 2604 176 2615 210
rect 2649 176 2661 210
rect 2604 120 2661 176
rect 2604 86 2615 120
rect 2649 86 2661 120
rect 2604 74 2661 86
rect 1536 48 1548 74
rect 1490 36 1548 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 464 86 476
rect 116 580 186 592
rect 116 546 139 580
rect 173 546 186 580
rect 116 510 186 546
rect 116 476 139 510
rect 173 476 186 510
rect 116 464 186 476
rect 216 464 270 592
rect 300 580 508 592
rect 300 546 313 580
rect 347 546 387 580
rect 421 546 461 580
rect 495 546 508 580
rect 300 510 508 546
rect 300 476 313 510
rect 347 476 387 510
rect 421 476 461 510
rect 495 476 508 510
rect 300 464 508 476
rect 538 464 592 592
rect 622 575 706 592
rect 622 541 635 575
rect 669 541 706 575
rect 622 464 706 541
rect 736 580 795 592
rect 736 546 749 580
rect 783 546 795 580
rect 736 510 795 546
rect 736 476 749 510
rect 783 476 795 510
rect 736 464 795 476
rect 855 421 914 592
rect 855 387 867 421
rect 901 387 914 421
rect 855 368 914 387
rect 944 580 1004 592
rect 944 546 957 580
rect 991 546 1004 580
rect 944 368 1004 546
rect 1034 421 1093 592
rect 1034 387 1047 421
rect 1081 387 1093 421
rect 1034 368 1093 387
rect 1445 582 1504 594
rect 1445 548 1457 582
rect 1491 548 1504 582
rect 1445 545 1504 548
rect 1862 560 1963 592
rect 1862 547 1895 560
rect 1260 541 1313 545
rect 1153 516 1212 541
rect 1153 482 1165 516
rect 1199 482 1212 516
rect 1153 457 1212 482
rect 1242 528 1313 541
rect 1242 494 1266 528
rect 1300 494 1313 528
rect 1242 461 1313 494
rect 1343 461 1397 545
rect 1427 461 1522 545
rect 1552 523 1611 545
rect 1552 489 1565 523
rect 1599 489 1611 523
rect 1552 461 1611 489
rect 1665 535 1724 547
rect 1665 501 1677 535
rect 1711 501 1724 535
rect 1665 467 1724 501
rect 1242 457 1295 461
rect 1665 433 1677 467
rect 1711 433 1724 467
rect 1665 399 1724 433
rect 1665 365 1677 399
rect 1711 365 1724 399
rect 1665 347 1724 365
rect 1754 535 1814 547
rect 1754 501 1767 535
rect 1801 501 1814 535
rect 1754 464 1814 501
rect 1754 430 1767 464
rect 1801 430 1814 464
rect 1754 393 1814 430
rect 1754 359 1767 393
rect 1801 359 1814 393
rect 1754 347 1814 359
rect 1844 526 1895 547
rect 1929 526 1963 560
rect 1844 508 1963 526
rect 1993 508 2047 592
rect 2077 567 2162 592
rect 2077 533 2097 567
rect 2131 533 2162 567
rect 2077 508 2162 533
rect 2192 567 2252 592
rect 2192 533 2205 567
rect 2239 533 2252 567
rect 2192 508 2252 533
rect 2282 580 2369 592
rect 2282 546 2312 580
rect 2346 546 2369 580
rect 2282 508 2369 546
rect 1844 347 1897 508
rect 2300 470 2369 508
rect 2300 436 2312 470
rect 2346 436 2369 470
rect 2300 424 2369 436
rect 2399 580 2458 592
rect 2399 546 2412 580
rect 2446 546 2458 580
rect 2399 470 2458 546
rect 2399 436 2412 470
rect 2446 436 2458 470
rect 2399 424 2458 436
rect 2512 580 2571 592
rect 2512 546 2524 580
rect 2558 546 2571 580
rect 2512 497 2571 546
rect 2512 463 2524 497
rect 2558 463 2571 497
rect 2512 414 2571 463
rect 2512 380 2524 414
rect 2558 380 2571 414
rect 2512 368 2571 380
rect 2601 580 2660 592
rect 2601 546 2614 580
rect 2648 546 2660 580
rect 2601 497 2660 546
rect 2601 463 2614 497
rect 2648 463 2660 497
rect 2601 414 2660 463
rect 2601 380 2614 414
rect 2648 380 2660 414
rect 2601 368 2660 380
<< ndiffc >>
rect 39 113 73 147
rect 873 168 907 202
rect 125 113 159 147
rect 237 93 271 127
rect 470 119 504 153
rect 652 93 686 127
rect 757 96 791 130
rect 873 86 907 120
rect 959 93 993 127
rect 1046 176 1080 210
rect 1046 86 1080 120
rect 1158 145 1192 179
rect 1244 145 1278 179
rect 1502 48 1536 82
rect 1670 145 1704 179
rect 1897 95 1931 129
rect 2055 99 2089 133
rect 2218 99 2252 133
rect 2330 83 2364 117
rect 2417 112 2451 146
rect 2529 176 2563 210
rect 2529 86 2563 120
rect 2615 176 2649 210
rect 2615 86 2649 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 139 546 173 580
rect 139 476 173 510
rect 313 546 347 580
rect 387 546 421 580
rect 461 546 495 580
rect 313 476 347 510
rect 387 476 421 510
rect 461 476 495 510
rect 635 541 669 575
rect 749 546 783 580
rect 749 476 783 510
rect 867 387 901 421
rect 957 546 991 580
rect 1047 387 1081 421
rect 1457 548 1491 582
rect 1165 482 1199 516
rect 1266 494 1300 528
rect 1565 489 1599 523
rect 1677 501 1711 535
rect 1677 433 1711 467
rect 1677 365 1711 399
rect 1767 501 1801 535
rect 1767 430 1801 464
rect 1767 359 1801 393
rect 1895 526 1929 560
rect 2097 533 2131 567
rect 2205 533 2239 567
rect 2312 546 2346 580
rect 2312 436 2346 470
rect 2412 546 2446 580
rect 2412 436 2446 470
rect 2524 546 2558 580
rect 2524 463 2558 497
rect 2524 380 2558 414
rect 2614 546 2648 580
rect 2614 463 2648 497
rect 2614 380 2648 414
<< poly >>
rect 86 592 116 618
rect 186 592 216 618
rect 270 592 300 618
rect 508 592 538 618
rect 592 592 622 618
rect 706 592 736 618
rect 914 592 944 618
rect 1004 592 1034 618
rect 1108 615 1847 645
rect 86 449 116 464
rect 186 449 216 464
rect 270 449 300 464
rect 508 449 538 464
rect 592 449 622 464
rect 706 449 736 464
rect 83 367 119 449
rect 183 367 219 449
rect 267 445 303 449
rect 267 415 353 445
rect 505 432 541 449
rect 83 351 225 367
rect 83 337 107 351
rect 84 317 107 337
rect 141 317 175 351
rect 209 317 225 351
rect 84 301 225 317
rect 323 318 353 415
rect 407 416 541 432
rect 407 382 423 416
rect 457 382 491 416
rect 525 382 541 416
rect 407 366 541 382
rect 589 422 625 449
rect 703 432 739 449
rect 589 406 655 422
rect 589 372 605 406
rect 639 372 655 406
rect 703 416 823 432
rect 703 402 773 416
rect 589 338 655 372
rect 84 172 114 301
rect 323 288 384 318
rect 354 253 384 288
rect 479 302 545 318
rect 479 268 495 302
rect 529 268 545 302
rect 589 304 605 338
rect 639 304 655 338
rect 589 288 655 304
rect 716 382 773 402
rect 807 382 823 416
rect 716 366 823 382
rect 209 237 275 253
rect 209 203 225 237
rect 259 217 275 237
rect 354 237 420 253
rect 479 252 545 268
rect 259 203 312 217
rect 209 187 312 203
rect 354 203 370 237
rect 404 203 420 237
rect 354 187 420 203
rect 282 165 312 187
rect 360 165 390 187
rect 515 165 545 252
rect 593 165 623 288
rect 716 165 746 366
rect 914 353 944 368
rect 1004 353 1034 368
rect 911 318 947 353
rect 1001 326 1037 353
rect 794 302 948 318
rect 794 268 810 302
rect 844 268 878 302
rect 912 268 948 302
rect 794 252 948 268
rect 918 222 948 252
rect 990 310 1056 326
rect 990 276 1006 310
rect 1040 276 1056 310
rect 990 267 1056 276
rect 1108 267 1138 615
rect 1212 541 1242 567
rect 1310 560 1346 615
rect 1313 545 1343 560
rect 1397 545 1427 571
rect 1522 545 1552 571
rect 1724 547 1754 573
rect 1811 562 1847 615
rect 1963 592 1993 618
rect 2047 592 2077 618
rect 2162 592 2192 618
rect 2252 592 2282 618
rect 2369 592 2399 618
rect 2571 592 2601 618
rect 1814 547 1844 562
rect 1212 442 1242 457
rect 1209 375 1245 442
rect 1313 435 1343 461
rect 1397 446 1427 461
rect 1522 446 1552 461
rect 1180 359 1246 375
rect 1394 361 1430 446
rect 1519 429 1555 446
rect 1519 413 1633 429
rect 1519 379 1583 413
rect 1617 379 1633 413
rect 1519 363 1633 379
rect 1180 325 1196 359
rect 1230 345 1246 359
rect 1367 345 1470 361
rect 1230 325 1319 345
rect 1180 315 1319 325
rect 1180 309 1246 315
rect 990 237 1233 267
rect 1005 222 1035 237
rect 84 62 114 88
rect 282 55 312 81
rect 360 55 390 81
rect 515 55 545 81
rect 593 55 623 81
rect 716 55 746 81
rect 1203 202 1233 237
rect 1289 202 1319 315
rect 1367 311 1420 345
rect 1454 311 1470 345
rect 1367 295 1470 311
rect 1367 202 1397 295
rect 1519 247 1549 363
rect 1963 493 1993 508
rect 2047 493 2077 508
rect 2162 493 2192 508
rect 2252 493 2282 508
rect 1960 476 1996 493
rect 1929 460 1996 476
rect 1929 426 1945 460
rect 1979 426 1996 460
rect 1929 410 1996 426
rect 2044 368 2080 493
rect 2159 430 2195 493
rect 1724 332 1754 347
rect 1814 332 1844 347
rect 2033 338 2080 368
rect 2128 414 2195 430
rect 2128 380 2144 414
rect 2178 380 2195 414
rect 2128 364 2195 380
rect 2249 398 2285 493
rect 2369 409 2399 424
rect 2366 398 2402 409
rect 2249 368 2402 398
rect 1721 319 1757 332
rect 1633 315 1757 319
rect 1597 299 1757 315
rect 1811 302 1955 332
rect 1597 265 1613 299
rect 1647 289 1757 299
rect 1647 265 1663 289
rect 1597 249 1663 265
rect 1445 217 1549 247
rect 1445 202 1475 217
rect 1629 202 1659 249
rect 1817 247 1883 254
rect 1715 238 1883 247
rect 1715 217 1833 238
rect 1715 202 1745 217
rect 1817 204 1833 217
rect 1867 204 1883 238
rect 1203 92 1233 118
rect 1289 92 1319 118
rect 1367 92 1397 118
rect 1445 92 1475 118
rect 918 48 948 74
rect 1005 48 1035 74
rect 1817 188 1883 204
rect 1925 224 1955 302
rect 1997 322 2063 338
rect 1997 288 2013 322
rect 2047 288 2063 322
rect 2128 290 2158 364
rect 1997 272 2063 288
rect 1925 194 1972 224
rect 1942 158 1972 194
rect 2014 158 2044 272
rect 2105 260 2158 290
rect 2249 270 2279 368
rect 2571 353 2601 368
rect 2568 326 2604 353
rect 2448 310 2604 326
rect 2448 276 2464 310
rect 2498 276 2532 310
rect 2566 276 2604 310
rect 2105 158 2135 260
rect 2213 254 2406 270
rect 2448 260 2604 276
rect 2213 220 2229 254
rect 2263 240 2406 254
rect 2263 220 2279 240
rect 2213 218 2279 220
rect 2177 188 2279 218
rect 2177 158 2207 188
rect 2376 184 2406 240
rect 2574 222 2604 260
rect 1629 48 1659 74
rect 1715 48 1745 74
rect 1942 48 1972 74
rect 2014 48 2044 74
rect 2105 48 2135 74
rect 2177 48 2207 74
rect 2376 48 2406 74
rect 2574 48 2604 74
<< polycont >>
rect 107 317 141 351
rect 175 317 209 351
rect 423 382 457 416
rect 491 382 525 416
rect 605 372 639 406
rect 495 268 529 302
rect 605 304 639 338
rect 773 382 807 416
rect 225 203 259 237
rect 370 203 404 237
rect 810 268 844 302
rect 878 268 912 302
rect 1006 276 1040 310
rect 1583 379 1617 413
rect 1196 325 1230 359
rect 1420 311 1454 345
rect 1945 426 1979 460
rect 2144 380 2178 414
rect 1613 265 1647 299
rect 1833 204 1867 238
rect 2013 288 2047 322
rect 2464 276 2498 310
rect 2532 276 2566 310
rect 2229 220 2263 254
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 435 89 476
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 510 189 546
rect 123 476 139 510
rect 173 476 189 510
rect 123 469 189 476
rect 297 580 511 596
rect 297 546 313 580
rect 347 546 387 580
rect 421 546 461 580
rect 495 546 511 580
rect 297 510 511 546
rect 619 575 685 649
rect 619 541 635 575
rect 669 541 685 575
rect 619 537 685 541
rect 733 580 799 596
rect 733 546 749 580
rect 783 546 799 580
rect 941 580 1007 649
rect 941 546 957 580
rect 991 546 1007 580
rect 1441 582 1508 649
rect 1441 548 1457 582
rect 1491 548 1508 582
rect 297 476 313 510
rect 347 476 387 510
rect 421 476 461 510
rect 495 503 511 510
rect 733 512 799 546
rect 1165 516 1215 545
rect 733 510 1165 512
rect 733 503 749 510
rect 495 476 749 503
rect 783 482 1165 510
rect 1199 482 1215 516
rect 783 478 1215 482
rect 783 476 799 478
rect 297 469 799 476
rect 689 466 799 469
rect 23 416 541 435
rect 23 401 423 416
rect 23 253 57 401
rect 407 382 423 401
rect 457 382 491 416
rect 525 382 541 416
rect 91 351 359 367
rect 407 366 541 382
rect 589 406 655 430
rect 589 372 605 406
rect 639 372 655 406
rect 91 317 107 351
rect 141 317 175 351
rect 209 332 359 351
rect 589 338 655 372
rect 209 317 545 332
rect 91 302 545 317
rect 91 298 495 302
rect 479 268 495 298
rect 529 268 545 302
rect 589 304 605 338
rect 639 304 655 338
rect 589 288 655 304
rect 23 237 275 253
rect 23 210 225 237
rect 23 147 73 210
rect 209 203 225 210
rect 259 203 275 237
rect 209 187 275 203
rect 313 237 420 253
rect 479 252 545 268
rect 313 203 370 237
rect 404 203 420 237
rect 689 218 723 466
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 807 382 833 390
rect 757 366 833 382
rect 867 421 917 444
rect 901 398 917 421
rect 1031 421 1124 444
rect 901 387 996 398
rect 867 364 996 387
rect 1031 387 1047 421
rect 1081 387 1124 421
rect 1165 443 1215 478
rect 1250 528 1376 545
rect 1441 532 1508 548
rect 1250 494 1266 528
rect 1300 498 1376 528
rect 1549 523 1615 549
rect 1549 498 1565 523
rect 1300 494 1565 498
rect 1250 489 1565 494
rect 1599 489 1615 523
rect 1250 477 1615 489
rect 1342 464 1615 477
rect 1677 535 1711 649
rect 1858 560 2063 576
rect 1677 467 1711 501
rect 1165 409 1308 443
rect 1031 375 1124 387
rect 1031 364 1240 375
rect 962 326 996 364
rect 1090 359 1240 364
rect 793 302 928 318
rect 793 268 810 302
rect 844 268 878 302
rect 912 268 928 302
rect 793 252 928 268
rect 962 310 1056 326
rect 962 276 1006 310
rect 1040 276 1056 310
rect 962 260 1056 276
rect 1090 325 1196 359
rect 1230 325 1240 359
rect 1090 309 1240 325
rect 793 236 839 252
rect 962 218 996 260
rect 1090 226 1124 309
rect 1274 274 1308 409
rect 23 113 39 147
rect 23 84 73 113
rect 109 147 175 176
rect 313 162 420 203
rect 454 184 723 218
rect 873 202 996 218
rect 109 113 125 147
rect 159 113 175 147
rect 454 153 520 184
rect 109 17 175 113
rect 221 127 287 128
rect 221 93 237 127
rect 271 93 287 127
rect 454 119 470 153
rect 504 119 520 153
rect 907 184 996 202
rect 1030 210 1124 226
rect 618 127 721 143
rect 221 85 287 93
rect 618 93 652 127
rect 686 93 721 127
rect 618 85 721 93
rect 221 51 721 85
rect 757 130 791 150
rect 757 17 791 96
rect 873 120 907 168
rect 1030 176 1046 210
rect 1080 176 1124 210
rect 873 70 907 86
rect 943 127 993 150
rect 943 93 959 127
rect 943 17 993 93
rect 1030 120 1124 176
rect 1030 86 1046 120
rect 1080 86 1124 120
rect 1158 240 1308 274
rect 1158 179 1192 240
rect 1342 206 1376 464
rect 1158 119 1192 145
rect 1228 179 1376 206
rect 1410 345 1465 361
rect 1410 311 1420 345
rect 1454 311 1465 345
rect 1410 218 1465 311
rect 1499 315 1533 464
rect 1567 424 1633 430
rect 1601 413 1633 424
rect 1567 379 1583 390
rect 1617 379 1633 413
rect 1567 363 1633 379
rect 1677 399 1711 433
rect 1677 349 1711 365
rect 1745 535 1801 551
rect 1745 501 1767 535
rect 1858 526 1895 560
rect 1929 526 2063 560
rect 1858 510 2063 526
rect 1745 464 1801 501
rect 1745 430 1767 464
rect 1745 393 1801 430
rect 1745 359 1767 393
rect 1745 343 1801 359
rect 1849 460 1995 476
rect 1849 426 1945 460
rect 1979 426 1995 460
rect 1849 425 1995 426
rect 1499 299 1663 315
rect 1499 265 1613 299
rect 1647 265 1663 299
rect 1499 252 1663 265
rect 1745 218 1779 343
rect 1849 254 1883 425
rect 2029 391 2063 510
rect 2097 567 2147 649
rect 2131 533 2147 567
rect 2097 504 2147 533
rect 2189 567 2262 596
rect 2189 533 2205 567
rect 2239 533 2262 567
rect 2189 504 2262 533
rect 1410 184 1779 218
rect 1813 238 1883 254
rect 1813 204 1833 238
rect 1867 204 1883 238
rect 1813 188 1883 204
rect 1917 357 2063 391
rect 2128 424 2194 430
rect 2128 390 2143 424
rect 2177 414 2194 424
rect 2128 380 2144 390
rect 2178 380 2194 414
rect 2128 364 2194 380
rect 1917 253 1951 357
rect 2228 323 2262 504
rect 2296 580 2362 649
rect 2296 546 2312 580
rect 2346 546 2362 580
rect 2296 470 2362 546
rect 2296 436 2312 470
rect 2346 436 2362 470
rect 2296 420 2362 436
rect 2396 580 2462 596
rect 2396 546 2412 580
rect 2446 546 2462 580
rect 2396 470 2462 546
rect 2396 436 2412 470
rect 2446 436 2462 470
rect 2396 420 2462 436
rect 2417 326 2462 420
rect 2508 580 2574 649
rect 2508 546 2524 580
rect 2558 546 2574 580
rect 2508 497 2574 546
rect 2508 463 2524 497
rect 2558 463 2574 497
rect 2508 414 2574 463
rect 2508 380 2524 414
rect 2558 380 2574 414
rect 2508 364 2574 380
rect 2614 580 2665 596
rect 2648 546 2665 580
rect 2614 497 2665 546
rect 2648 463 2665 497
rect 2614 414 2665 463
rect 2648 380 2665 414
rect 1997 322 2347 323
rect 1997 288 2013 322
rect 2047 289 2347 322
rect 2047 288 2063 289
rect 1997 287 2063 288
rect 2213 254 2279 255
rect 2213 253 2229 254
rect 1917 220 2229 253
rect 2263 220 2279 254
rect 1917 219 2279 220
rect 1228 145 1244 179
rect 1278 172 1376 179
rect 1654 179 1731 184
rect 1278 145 1294 172
rect 1228 119 1294 145
rect 1030 85 1124 86
rect 1410 116 1620 150
rect 1654 145 1670 179
rect 1704 145 1731 179
rect 1654 119 1731 145
rect 1410 85 1444 116
rect 1030 51 1444 85
rect 1586 85 1620 116
rect 1813 85 1847 188
rect 1917 154 1951 219
rect 2313 185 2347 289
rect 1486 48 1502 82
rect 1536 48 1552 82
rect 1586 51 1847 85
rect 1881 129 1951 154
rect 1881 95 1897 129
rect 1931 95 1951 129
rect 1881 70 1951 95
rect 2039 133 2105 162
rect 2039 99 2055 133
rect 2089 99 2105 133
rect 1486 17 1552 48
rect 2039 17 2105 99
rect 2202 151 2347 185
rect 2417 310 2574 326
rect 2417 276 2464 310
rect 2498 276 2532 310
rect 2566 276 2574 310
rect 2417 260 2574 276
rect 2202 133 2268 151
rect 2202 99 2218 133
rect 2252 99 2268 133
rect 2417 146 2467 260
rect 2614 226 2665 380
rect 2202 70 2268 99
rect 2314 83 2330 117
rect 2364 83 2381 117
rect 2314 17 2381 83
rect 2451 112 2467 146
rect 2417 70 2467 112
rect 2513 210 2563 226
rect 2513 176 2529 210
rect 2513 120 2563 176
rect 2513 86 2529 120
rect 2513 17 2563 86
rect 2599 210 2665 226
rect 2599 176 2615 210
rect 2649 176 2665 210
rect 2599 120 2665 176
rect 2599 86 2615 120
rect 2649 86 2665 120
rect 2599 70 2665 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1567 413 1601 424
rect 1567 390 1583 413
rect 1583 390 1601 413
rect 2143 414 2177 424
rect 2143 390 2144 414
rect 2144 390 2177 414
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfrtp_1
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel nbase s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel metal1 s 2143 390 2177 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew
flabel corelocali s 2623 94 2657 128 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 10 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew
flabel corelocali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew
flabel corelocali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2688 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 235530
string GDS_START 215032
<< end >>
