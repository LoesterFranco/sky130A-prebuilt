magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 55 427 89 527
rect 139 409 173 493
rect 207 443 273 527
rect 307 409 341 493
rect 375 443 441 527
rect 941 447 1007 527
rect 1783 455 1849 527
rect 139 291 341 409
rect 139 288 284 291
rect 221 185 284 288
rect 119 166 307 185
rect 119 132 321 166
rect 35 17 69 109
rect 119 70 153 132
rect 187 17 253 93
rect 287 70 321 132
rect 371 17 405 105
rect 576 199 703 265
rect 990 17 1024 177
rect 1541 289 1657 323
rect 1541 199 1575 289
rect 1705 215 1787 265
rect 1799 17 1833 113
rect 0 -17 2024 17
<< obsli1 >>
rect 475 447 783 481
rect 826 447 907 481
rect 1074 455 1693 489
rect 475 409 509 447
rect 873 413 907 447
rect 1074 413 1108 455
rect 375 375 509 409
rect 578 379 839 413
rect 873 379 1108 413
rect 375 265 409 375
rect 474 307 771 341
rect 364 193 409 265
rect 375 173 409 193
rect 375 139 473 173
rect 439 85 473 139
rect 508 119 542 307
rect 737 265 771 307
rect 805 339 839 379
rect 805 323 911 339
rect 805 305 877 323
rect 854 289 877 305
rect 854 275 911 289
rect 737 199 811 265
rect 598 131 820 165
rect 682 85 752 91
rect 439 51 752 85
rect 786 85 820 131
rect 854 119 888 275
rect 945 241 979 379
rect 1025 289 1108 343
rect 922 210 979 241
rect 922 209 978 210
rect 922 208 976 209
rect 922 207 973 208
rect 922 85 956 207
rect 1060 187 1108 289
rect 786 51 956 85
rect 1060 153 1061 187
rect 1095 153 1108 187
rect 1060 83 1108 153
rect 1143 119 1177 421
rect 1215 178 1249 455
rect 1883 421 1935 493
rect 1283 323 1366 409
rect 1473 387 1935 421
rect 1283 289 1337 323
rect 1371 289 1439 323
rect 1286 199 1371 254
rect 1328 187 1371 199
rect 1215 165 1255 178
rect 1215 144 1294 165
rect 1221 131 1294 144
rect 1143 85 1153 119
rect 1187 85 1226 97
rect 1143 53 1226 85
rect 1260 64 1294 131
rect 1328 153 1337 187
rect 1328 126 1371 153
rect 1405 85 1439 289
rect 1473 119 1507 387
rect 1838 375 1935 387
rect 1691 299 1855 341
rect 1821 265 1855 299
rect 1609 189 1671 255
rect 1821 199 1867 265
rect 1609 187 1650 189
rect 1609 153 1613 187
rect 1647 153 1650 187
rect 1821 181 1855 199
rect 1609 146 1650 153
rect 1707 150 1855 181
rect 1699 147 1855 150
rect 1699 119 1757 147
rect 1541 85 1634 93
rect 1405 51 1634 85
rect 1699 85 1705 119
rect 1739 85 1757 119
rect 1901 117 1935 375
rect 1699 59 1757 85
rect 1883 51 1935 117
<< obsli1c >>
rect 877 289 911 323
rect 1061 153 1095 187
rect 1337 289 1371 323
rect 1153 85 1187 119
rect 1337 153 1371 187
rect 1613 153 1647 187
rect 1705 85 1739 119
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< obsm1 >>
rect 865 323 923 329
rect 865 289 877 323
rect 911 320 923 323
rect 1325 323 1383 329
rect 1325 320 1337 323
rect 911 292 1337 320
rect 911 289 923 292
rect 865 283 923 289
rect 1325 289 1337 292
rect 1371 289 1383 323
rect 1325 283 1383 289
rect 1049 187 1107 193
rect 1049 153 1061 187
rect 1095 184 1107 187
rect 1325 187 1383 193
rect 1325 184 1337 187
rect 1095 156 1337 184
rect 1095 153 1107 156
rect 1049 147 1107 153
rect 1325 153 1337 156
rect 1371 184 1383 187
rect 1601 187 1659 193
rect 1601 184 1613 187
rect 1371 156 1613 184
rect 1371 153 1383 156
rect 1325 147 1383 153
rect 1601 153 1613 156
rect 1647 153 1659 187
rect 1601 147 1659 153
rect 1141 119 1199 125
rect 1141 85 1153 119
rect 1187 116 1199 119
rect 1693 119 1751 125
rect 1693 116 1705 119
rect 1187 88 1705 116
rect 1187 85 1199 88
rect 1141 79 1199 85
rect 1693 85 1705 88
rect 1739 85 1751 119
rect 1693 79 1751 85
<< labels >>
rlabel locali s 1705 215 1787 265 6 A
port 1 nsew signal input
rlabel locali s 1541 289 1657 323 6 B
port 2 nsew signal input
rlabel locali s 1541 199 1575 289 6 B
port 2 nsew signal input
rlabel locali s 576 199 703 265 6 C
port 3 nsew signal input
rlabel locali s 307 409 341 493 6 X
port 4 nsew signal output
rlabel locali s 287 70 321 132 6 X
port 4 nsew signal output
rlabel locali s 221 185 284 288 6 X
port 4 nsew signal output
rlabel locali s 139 409 173 493 6 X
port 4 nsew signal output
rlabel locali s 139 291 341 409 6 X
port 4 nsew signal output
rlabel locali s 139 288 284 291 6 X
port 4 nsew signal output
rlabel locali s 119 166 307 185 6 X
port 4 nsew signal output
rlabel locali s 119 132 321 166 6 X
port 4 nsew signal output
rlabel locali s 119 70 153 132 6 X
port 4 nsew signal output
rlabel locali s 1799 17 1833 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 990 17 1024 177 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 371 17 405 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 187 17 253 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 35 17 69 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1783 455 1849 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 941 447 1007 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 375 443 441 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 207 443 273 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 55 427 89 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 698948
string GDS_START 685650
<< end >>
