magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1012 561
rect 103 427 169 527
rect 291 451 370 527
rect 18 197 66 325
rect 350 153 425 219
rect 671 427 705 527
rect 859 314 893 527
rect 938 334 995 491
rect 103 17 169 93
rect 961 149 995 334
rect 291 17 357 93
rect 653 17 719 106
rect 859 17 893 143
rect 938 83 995 149
rect 0 -17 1012 17
<< obsli1 >>
rect 35 393 69 493
rect 203 417 237 493
rect 462 451 637 485
rect 203 393 569 417
rect 35 359 156 393
rect 122 292 156 359
rect 196 383 569 393
rect 196 365 237 383
rect 122 226 162 292
rect 122 161 156 226
rect 35 127 156 161
rect 196 182 230 365
rect 264 305 467 339
rect 264 248 298 305
rect 410 271 467 305
rect 501 315 569 383
rect 196 148 237 182
rect 501 207 535 315
rect 603 265 637 451
rect 767 373 825 487
rect 684 307 825 373
rect 603 233 756 265
rect 35 69 69 127
rect 203 69 237 148
rect 459 141 535 207
rect 574 199 756 233
rect 574 107 608 199
rect 790 149 825 307
rect 476 73 608 107
rect 767 83 825 149
<< metal1 >>
rect 0 496 1012 592
rect 0 -48 1012 48
<< labels >>
rlabel locali s 350 153 425 219 6 D
port 1 nsew signal input
rlabel locali s 961 149 995 334 6 Q
port 2 nsew signal output
rlabel locali s 938 334 995 491 6 Q
port 2 nsew signal output
rlabel locali s 938 83 995 149 6 Q
port 2 nsew signal output
rlabel locali s 18 197 66 325 6 SLEEP_B
port 3 nsew clock input
rlabel locali s 859 17 893 143 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 653 17 719 106 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 291 17 357 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 1012 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 859 314 893 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 671 427 705 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 291 451 370 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 1012 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1012 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2321054
string GDS_START 2312122
<< end >>
