magic
tech sky130A
magscale 1 2
timestamp 1604502710
<< nwell >>
rect -38 332 326 704
<< pwell >>
rect 0 0 288 49
<< scpmos >>
rect 81 424 117 592
rect 171 424 207 592
<< nmoslvt >>
rect 98 74 128 158
<< ndiff >>
rect 27 127 98 158
rect 27 93 39 127
rect 73 93 98 127
rect 27 74 98 93
rect 128 132 178 158
rect 128 120 261 132
rect 128 86 139 120
rect 173 86 215 120
rect 249 86 261 120
rect 128 74 261 86
<< pdiff >>
rect 27 580 81 592
rect 27 546 37 580
rect 71 546 81 580
rect 27 470 81 546
rect 27 436 37 470
rect 71 436 81 470
rect 27 424 81 436
rect 117 575 171 592
rect 117 541 127 575
rect 161 541 171 575
rect 117 470 171 541
rect 117 436 127 470
rect 161 436 171 470
rect 117 424 171 436
rect 207 575 261 592
rect 207 541 217 575
rect 251 541 261 575
rect 207 424 261 541
<< ndiffc >>
rect 39 93 73 127
rect 139 86 173 120
rect 215 86 249 120
<< pdiffc >>
rect 37 546 71 580
rect 37 436 71 470
rect 127 541 161 575
rect 127 436 161 470
rect 217 541 251 575
<< poly >>
rect 81 592 117 618
rect 171 592 207 618
rect 81 386 117 424
rect 171 386 207 424
rect 81 370 207 386
rect 81 336 101 370
rect 135 336 207 370
rect 81 302 207 336
rect 81 268 101 302
rect 135 268 207 302
rect 81 234 207 268
rect 81 200 101 234
rect 135 200 207 234
rect 81 184 207 200
rect 98 158 128 184
rect 98 48 128 74
<< polycont >>
rect 101 336 135 370
rect 101 268 135 302
rect 101 200 135 234
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 21 580 71 649
rect 21 546 37 580
rect 21 470 71 546
rect 21 436 37 470
rect 21 420 71 436
rect 111 575 167 591
rect 111 541 127 575
rect 161 541 167 575
rect 111 486 167 541
rect 201 575 267 649
rect 201 541 217 575
rect 251 541 267 575
rect 201 520 267 541
rect 111 470 265 486
rect 111 436 127 470
rect 161 436 265 470
rect 111 420 265 436
rect 85 370 151 386
rect 85 356 101 370
rect 25 336 101 356
rect 135 336 151 370
rect 25 302 151 336
rect 25 268 101 302
rect 135 268 151 302
rect 25 236 151 268
rect 85 234 151 236
rect 85 200 101 234
rect 135 200 151 234
rect 85 184 151 200
rect 23 127 89 150
rect 217 136 265 420
rect 23 93 39 127
rect 73 93 89 127
rect 23 17 89 93
rect 123 120 265 136
rect 123 86 139 120
rect 173 86 215 120
rect 249 86 265 120
rect 123 70 265 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 683 288 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 0 617 288 649
rect 0 17 288 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -49 288 -17
<< labels >>
flabel pwell s 0 0 288 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 288 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 0 0 0 4 clkinv_1
flabel metal1 s 0 617 288 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 288 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 94 257 128 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 223 242 257 276 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 6 nsew
flabel corelocali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 288 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string GDS_END 2581942
string GDS_START 2578006
<< end >>
