magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 391 455 457 596
rect 321 390 457 455
rect 89 288 263 356
rect 321 226 355 390
rect 389 260 455 356
rect 321 192 457 226
rect 391 70 457 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 21 549 178 615
rect 21 402 176 549
rect 217 404 283 649
rect 21 212 55 402
rect 21 82 188 212
rect 227 17 284 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 389 260 455 356 6 A
port 1 nsew signal input
rlabel locali s 89 288 263 356 6 TE
port 2 nsew signal input
rlabel locali s 391 455 457 596 6 Z
port 3 nsew signal output
rlabel locali s 391 70 457 192 6 Z
port 3 nsew signal output
rlabel locali s 321 390 457 455 6 Z
port 3 nsew signal output
rlabel locali s 321 226 355 390 6 Z
port 3 nsew signal output
rlabel locali s 321 192 457 226 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 617 480 715 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2096046
string GDS_START 2091050
<< end >>
