magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scnmos >>
rect 121 74 151 222
rect 207 74 237 222
rect 369 74 399 222
rect 441 74 471 222
rect 549 74 579 222
rect 657 74 687 222
<< pmoshvt >>
rect 88 368 118 592
rect 178 368 208 592
rect 372 392 402 592
rect 480 392 510 592
rect 570 392 600 592
rect 654 392 684 592
<< ndiff >>
rect 68 136 121 222
rect 68 102 76 136
rect 110 102 121 136
rect 68 74 121 102
rect 151 210 207 222
rect 151 176 162 210
rect 196 176 207 210
rect 151 120 207 176
rect 151 86 162 120
rect 196 86 207 120
rect 151 74 207 86
rect 237 127 369 222
rect 237 93 248 127
rect 282 93 324 127
rect 358 93 369 127
rect 237 74 369 93
rect 399 74 441 222
rect 471 202 549 222
rect 471 168 486 202
rect 520 168 549 202
rect 471 120 549 168
rect 471 86 486 120
rect 520 86 549 120
rect 471 74 549 86
rect 579 127 657 222
rect 579 93 601 127
rect 635 93 657 127
rect 579 74 657 93
rect 687 210 740 222
rect 687 176 698 210
rect 732 176 740 210
rect 687 120 740 176
rect 687 86 698 120
rect 732 86 740 120
rect 687 74 740 86
<< pdiff >>
rect 33 580 88 592
rect 33 546 41 580
rect 75 546 88 580
rect 33 497 88 546
rect 33 463 41 497
rect 75 463 88 497
rect 33 414 88 463
rect 33 380 41 414
rect 75 380 88 414
rect 33 368 88 380
rect 118 580 178 592
rect 118 546 131 580
rect 165 546 178 580
rect 118 497 178 546
rect 118 463 131 497
rect 165 463 178 497
rect 118 414 178 463
rect 118 380 131 414
rect 165 380 178 414
rect 118 368 178 380
rect 208 580 263 592
rect 208 546 221 580
rect 255 546 263 580
rect 208 508 263 546
rect 208 474 221 508
rect 255 474 263 508
rect 208 368 263 474
rect 317 580 372 592
rect 317 546 325 580
rect 359 546 372 580
rect 317 508 372 546
rect 317 474 325 508
rect 359 474 372 508
rect 317 392 372 474
rect 402 578 480 592
rect 402 544 419 578
rect 453 544 480 578
rect 402 392 480 544
rect 510 580 570 592
rect 510 546 523 580
rect 557 546 570 580
rect 510 508 570 546
rect 510 474 523 508
rect 557 474 570 508
rect 510 392 570 474
rect 600 392 654 592
rect 684 580 739 592
rect 684 546 697 580
rect 731 546 739 580
rect 684 510 739 546
rect 684 476 697 510
rect 731 476 739 510
rect 684 440 739 476
rect 684 406 697 440
rect 731 406 739 440
rect 684 392 739 406
<< ndiffc >>
rect 76 102 110 136
rect 162 176 196 210
rect 162 86 196 120
rect 248 93 282 127
rect 324 93 358 127
rect 486 168 520 202
rect 486 86 520 120
rect 601 93 635 127
rect 698 176 732 210
rect 698 86 732 120
<< pdiffc >>
rect 41 546 75 580
rect 41 463 75 497
rect 41 380 75 414
rect 131 546 165 580
rect 131 463 165 497
rect 131 380 165 414
rect 221 546 255 580
rect 221 474 255 508
rect 325 546 359 580
rect 325 474 359 508
rect 419 544 453 578
rect 523 546 557 580
rect 523 474 557 508
rect 697 546 731 580
rect 697 476 731 510
rect 697 406 731 440
<< poly >>
rect 88 592 118 618
rect 178 592 208 618
rect 372 592 402 618
rect 480 592 510 618
rect 570 592 600 618
rect 654 592 684 618
rect 372 377 402 392
rect 480 377 510 392
rect 570 377 600 392
rect 654 377 684 392
rect 88 353 118 368
rect 178 353 208 368
rect 85 300 121 353
rect 175 336 211 353
rect 369 346 405 377
rect 477 346 513 377
rect 175 320 267 336
rect 175 300 217 320
rect 85 286 217 300
rect 251 286 267 320
rect 369 318 399 346
rect 477 318 507 346
rect 567 318 603 377
rect 651 356 687 377
rect 651 346 747 356
rect 657 340 747 346
rect 85 270 267 286
rect 309 302 399 318
rect 121 222 151 270
rect 207 222 237 270
rect 309 268 325 302
rect 359 268 399 302
rect 309 252 399 268
rect 369 222 399 252
rect 441 302 507 318
rect 441 268 457 302
rect 491 268 507 302
rect 441 252 507 268
rect 549 302 615 318
rect 549 268 565 302
rect 599 268 615 302
rect 549 252 615 268
rect 657 306 697 340
rect 731 306 747 340
rect 657 290 747 306
rect 441 222 471 252
rect 549 222 579 252
rect 657 222 687 290
rect 121 48 151 74
rect 207 48 237 74
rect 369 48 399 74
rect 441 48 471 74
rect 549 48 579 74
rect 657 48 687 74
<< polycont >>
rect 217 286 251 320
rect 325 268 359 302
rect 457 268 491 302
rect 565 268 599 302
rect 697 306 731 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 580 75 649
rect 25 546 41 580
rect 25 497 75 546
rect 25 463 41 497
rect 25 414 75 463
rect 25 380 41 414
rect 25 364 75 380
rect 115 580 167 596
rect 115 546 131 580
rect 165 546 167 580
rect 115 497 167 546
rect 115 463 131 497
rect 165 463 167 497
rect 115 414 167 463
rect 205 580 271 649
rect 205 546 221 580
rect 255 546 271 580
rect 205 508 271 546
rect 205 474 221 508
rect 255 474 271 508
rect 205 458 271 474
rect 309 580 375 596
rect 309 546 325 580
rect 359 546 375 580
rect 309 508 375 546
rect 415 578 473 649
rect 415 544 419 578
rect 453 544 473 578
rect 415 526 473 544
rect 507 580 573 596
rect 507 546 523 580
rect 557 546 573 580
rect 309 474 325 508
rect 359 492 375 508
rect 507 508 573 546
rect 507 492 523 508
rect 359 474 523 492
rect 557 474 573 508
rect 309 458 573 474
rect 681 580 747 596
rect 681 546 697 580
rect 731 546 747 580
rect 681 510 747 546
rect 681 476 697 510
rect 731 476 747 510
rect 681 440 747 476
rect 681 424 697 440
rect 115 380 131 414
rect 165 380 167 414
rect 115 236 167 380
rect 233 406 697 424
rect 731 406 747 440
rect 233 390 747 406
rect 233 336 267 390
rect 201 320 267 336
rect 201 286 217 320
rect 251 286 267 320
rect 201 270 267 286
rect 115 210 196 236
rect 115 202 162 210
rect 233 218 267 270
rect 309 302 375 356
rect 309 268 325 302
rect 359 268 375 302
rect 309 252 375 268
rect 409 302 507 356
rect 409 268 457 302
rect 491 268 507 302
rect 409 252 507 268
rect 549 302 647 356
rect 549 268 565 302
rect 599 268 647 302
rect 681 340 747 356
rect 681 306 697 340
rect 731 306 747 340
rect 681 290 747 306
rect 549 252 647 268
rect 698 218 748 226
rect 233 210 748 218
rect 233 202 698 210
rect 233 184 486 202
rect 60 136 126 168
rect 60 102 76 136
rect 110 102 126 136
rect 60 17 126 102
rect 162 120 196 176
rect 466 168 486 184
rect 520 184 698 202
rect 520 168 540 184
rect 162 70 196 86
rect 232 127 374 150
rect 232 93 248 127
rect 282 93 324 127
rect 358 93 374 127
rect 232 70 374 93
rect 466 120 540 168
rect 732 176 748 210
rect 466 86 486 120
rect 520 86 540 120
rect 466 70 540 86
rect 574 127 662 150
rect 574 93 601 127
rect 635 93 662 127
rect 574 70 662 93
rect 698 120 748 176
rect 732 86 748 120
rect 698 70 748 86
rect 232 17 266 70
rect 574 17 608 70
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a211o_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 4 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel corelocali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3939118
string GDS_START 3931714
<< end >>
