magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 21 271 111 353
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 118 462 177 649
rect 20 428 86 445
rect 20 387 179 428
rect 145 321 179 387
rect 213 424 276 615
rect 420 462 479 649
rect 213 390 223 424
rect 257 390 276 424
rect 213 367 276 390
rect 310 428 374 445
rect 513 432 573 615
rect 717 462 776 649
rect 310 379 467 428
rect 242 321 276 367
rect 433 321 467 379
rect 501 424 573 432
rect 501 390 511 424
rect 545 390 573 424
rect 501 367 573 390
rect 614 428 680 445
rect 810 432 870 615
rect 614 379 761 428
rect 539 321 573 367
rect 721 321 761 379
rect 795 424 870 432
rect 795 390 799 424
rect 833 390 870 424
rect 795 367 870 390
rect 145 255 208 321
rect 242 263 399 321
rect 145 229 179 255
rect 20 195 179 229
rect 242 215 276 263
rect 433 255 505 321
rect 539 263 687 321
rect 433 229 467 255
rect 20 140 79 195
rect 118 17 184 161
rect 218 51 276 215
rect 310 195 467 229
rect 539 215 573 263
rect 721 255 802 321
rect 721 229 755 255
rect 310 140 367 195
rect 406 17 472 161
rect 506 51 573 215
rect 612 195 755 229
rect 836 215 870 367
rect 612 140 655 195
rect 694 17 760 161
rect 794 51 870 215
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 223 390 257 424
rect 511 390 545 424
rect 799 390 833 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 193 464 842 498
rect 481 424 557 464
rect 481 390 511 424
rect 545 390 557 424
rect 481 384 557 390
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< obsm1 >>
rect 193 424 269 430
rect 193 390 223 424
rect 257 390 269 424
rect 193 384 269 390
rect 769 424 845 430
rect 769 390 799 424
rect 833 390 845 424
rect 769 384 845 390
<< labels >>
rlabel locali s 21 271 111 353 6 A
port 1 nsew signal input
rlabel metal1 s 481 384 557 464 6 X
port 2 nsew signal output
rlabel metal1 s 193 464 842 498 6 X
port 2 nsew signal output
rlabel metal1 s 0 -49 960 49 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 617 960 715 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2028950
string GDS_START 2020854
<< end >>
