magic
tech sky130A
magscale 1 2
timestamp 1604502705
<< nwell >>
rect -38 356 1574 704
rect -38 332 232 356
rect 871 351 1574 356
rect 1241 332 1574 351
<< pwell >>
rect 0 0 1536 49
<< scnmos >>
rect 84 74 114 222
rect 237 74 267 202
rect 315 74 345 202
rect 464 118 494 202
rect 559 139 589 223
rect 716 125 746 273
rect 914 119 944 267
rect 1014 119 1044 267
rect 1086 119 1116 267
rect 1336 92 1366 240
rect 1422 92 1452 240
<< pmoshvt >>
rect 86 368 116 592
rect 234 392 264 592
rect 318 392 348 592
rect 478 508 508 592
rect 562 508 592 592
rect 704 424 734 592
rect 910 419 940 587
rect 1011 387 1041 587
rect 1106 387 1136 587
rect 1330 368 1360 592
rect 1420 368 1450 592
<< ndiff >>
rect 27 146 84 222
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 202 164 222
rect 666 223 716 273
rect 509 202 559 223
rect 114 120 237 202
rect 114 86 125 120
rect 159 86 237 120
rect 114 74 237 86
rect 267 74 315 202
rect 345 174 464 202
rect 345 140 380 174
rect 414 140 464 174
rect 345 118 464 140
rect 494 139 559 202
rect 589 185 716 223
rect 589 151 600 185
rect 634 151 671 185
rect 705 151 716 185
rect 589 139 716 151
rect 494 118 544 139
rect 345 74 395 118
rect 666 125 716 139
rect 746 261 803 273
rect 746 227 757 261
rect 791 227 803 261
rect 746 171 803 227
rect 746 137 757 171
rect 791 137 803 171
rect 746 125 803 137
rect 857 239 914 267
rect 857 205 869 239
rect 903 205 914 239
rect 857 165 914 205
rect 857 131 869 165
rect 903 131 914 165
rect 857 119 914 131
rect 944 239 1014 267
rect 944 205 969 239
rect 1003 205 1014 239
rect 944 165 1014 205
rect 944 131 969 165
rect 1003 131 1014 165
rect 944 119 1014 131
rect 1044 119 1086 267
rect 1116 255 1173 267
rect 1116 221 1127 255
rect 1161 221 1173 255
rect 1116 165 1173 221
rect 1116 131 1127 165
rect 1161 131 1173 165
rect 1286 150 1336 240
rect 1116 119 1173 131
rect 1263 138 1336 150
rect 1263 104 1277 138
rect 1311 104 1336 138
rect 1263 92 1336 104
rect 1366 228 1422 240
rect 1366 194 1377 228
rect 1411 194 1422 228
rect 1366 138 1422 194
rect 1366 104 1377 138
rect 1411 104 1422 138
rect 1366 92 1422 104
rect 1452 228 1509 240
rect 1452 194 1463 228
rect 1497 194 1509 228
rect 1452 138 1509 194
rect 1452 104 1463 138
rect 1497 104 1509 138
rect 1452 92 1509 104
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 234 592
rect 116 546 159 580
rect 193 546 234 580
rect 116 494 234 546
rect 116 460 159 494
rect 193 460 234 494
rect 116 392 234 460
rect 264 392 318 592
rect 348 560 478 592
rect 348 526 361 560
rect 395 526 431 560
rect 465 526 478 560
rect 348 508 478 526
rect 508 508 562 592
rect 592 580 704 592
rect 592 546 626 580
rect 660 546 704 580
rect 592 508 704 546
rect 348 392 401 508
rect 116 368 169 392
rect 651 424 704 508
rect 734 580 793 592
rect 1265 587 1330 592
rect 734 546 747 580
rect 781 546 793 580
rect 734 470 793 546
rect 734 436 747 470
rect 781 436 793 470
rect 734 424 793 436
rect 847 575 910 587
rect 847 541 859 575
rect 893 541 910 575
rect 847 465 910 541
rect 847 431 859 465
rect 893 431 910 465
rect 847 419 910 431
rect 940 575 1011 587
rect 940 541 959 575
rect 993 541 1011 575
rect 940 465 1011 541
rect 940 431 959 465
rect 993 431 1011 465
rect 940 419 1011 431
rect 958 387 1011 419
rect 1041 579 1106 587
rect 1041 545 1059 579
rect 1093 545 1106 579
rect 1041 508 1106 545
rect 1041 474 1059 508
rect 1093 474 1106 508
rect 1041 436 1106 474
rect 1041 402 1059 436
rect 1093 402 1106 436
rect 1041 387 1106 402
rect 1136 579 1330 587
rect 1136 545 1150 579
rect 1184 545 1277 579
rect 1311 545 1330 579
rect 1136 508 1330 545
rect 1136 474 1150 508
rect 1184 474 1277 508
rect 1311 474 1330 508
rect 1136 440 1330 474
rect 1136 406 1150 440
rect 1184 406 1277 440
rect 1311 406 1330 440
rect 1136 387 1330 406
rect 1277 368 1330 387
rect 1360 580 1420 592
rect 1360 546 1373 580
rect 1407 546 1420 580
rect 1360 497 1420 546
rect 1360 463 1373 497
rect 1407 463 1420 497
rect 1360 414 1420 463
rect 1360 380 1373 414
rect 1407 380 1420 414
rect 1360 368 1420 380
rect 1450 580 1509 592
rect 1450 546 1463 580
rect 1497 546 1509 580
rect 1450 497 1509 546
rect 1450 463 1463 497
rect 1497 463 1509 497
rect 1450 414 1509 463
rect 1450 380 1463 414
rect 1497 380 1509 414
rect 1450 368 1509 380
<< ndiffc >>
rect 39 112 73 146
rect 125 86 159 120
rect 380 140 414 174
rect 600 151 634 185
rect 671 151 705 185
rect 757 227 791 261
rect 757 137 791 171
rect 869 205 903 239
rect 869 131 903 165
rect 969 205 1003 239
rect 969 131 1003 165
rect 1127 221 1161 255
rect 1127 131 1161 165
rect 1277 104 1311 138
rect 1377 194 1411 228
rect 1377 104 1411 138
rect 1463 194 1497 228
rect 1463 104 1497 138
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 159 546 193 580
rect 159 460 193 494
rect 361 526 395 560
rect 431 526 465 560
rect 626 546 660 580
rect 747 546 781 580
rect 747 436 781 470
rect 859 541 893 575
rect 859 431 893 465
rect 959 541 993 575
rect 959 431 993 465
rect 1059 545 1093 579
rect 1059 474 1093 508
rect 1059 402 1093 436
rect 1150 545 1184 579
rect 1277 545 1311 579
rect 1150 474 1184 508
rect 1277 474 1311 508
rect 1150 406 1184 440
rect 1277 406 1311 440
rect 1373 546 1407 580
rect 1373 463 1407 497
rect 1373 380 1407 414
rect 1463 546 1497 580
rect 1463 463 1497 497
rect 1463 380 1497 414
<< poly >>
rect 86 592 116 618
rect 234 592 264 618
rect 318 592 348 618
rect 478 592 508 618
rect 562 592 592 618
rect 704 592 734 618
rect 478 493 508 508
rect 562 493 592 508
rect 475 476 511 493
rect 445 460 511 476
rect 445 426 461 460
rect 495 426 511 460
rect 445 410 511 426
rect 559 425 595 493
rect 234 377 264 392
rect 318 377 348 392
rect 86 353 116 368
rect 231 356 267 377
rect 83 310 119 353
rect 201 340 267 356
rect 83 294 153 310
rect 83 260 103 294
rect 137 260 153 294
rect 201 306 217 340
rect 251 306 267 340
rect 315 368 351 377
rect 315 352 517 368
rect 315 338 467 352
rect 201 290 267 306
rect 451 318 467 338
rect 501 318 517 352
rect 451 302 517 318
rect 83 244 153 260
rect 84 222 114 244
rect 237 202 267 290
rect 315 274 409 290
rect 315 240 359 274
rect 393 240 409 274
rect 315 224 409 240
rect 315 202 345 224
rect 464 202 494 302
rect 559 223 589 425
rect 910 587 940 613
rect 1011 587 1041 613
rect 1106 587 1136 613
rect 1330 592 1360 618
rect 1420 592 1450 618
rect 704 409 734 424
rect 701 389 734 409
rect 910 404 940 419
rect 701 377 731 389
rect 631 361 731 377
rect 631 327 647 361
rect 681 341 731 361
rect 799 361 865 377
rect 799 341 815 361
rect 681 327 815 341
rect 849 327 865 361
rect 631 311 865 327
rect 907 355 943 404
rect 1011 372 1041 387
rect 1106 372 1136 387
rect 1008 355 1044 372
rect 907 339 1044 355
rect 716 273 746 311
rect 907 305 926 339
rect 960 305 994 339
rect 1028 305 1044 339
rect 1103 312 1139 372
rect 1330 353 1360 368
rect 1420 353 1450 368
rect 1327 322 1363 353
rect 1417 322 1453 353
rect 907 289 1044 305
rect 464 92 494 118
rect 559 117 589 139
rect 914 267 944 289
rect 1014 267 1044 289
rect 1086 282 1139 312
rect 1195 306 1453 322
rect 1086 267 1116 282
rect 1195 272 1211 306
rect 1245 274 1453 306
rect 1245 272 1261 274
rect 559 101 632 117
rect 84 48 114 74
rect 237 48 267 74
rect 315 48 345 74
rect 559 67 582 101
rect 616 67 632 101
rect 716 99 746 125
rect 1195 238 1261 272
rect 1336 240 1366 274
rect 1422 262 1453 274
rect 1422 240 1452 262
rect 1195 204 1211 238
rect 1245 204 1261 238
rect 1195 188 1261 204
rect 914 93 944 119
rect 1014 93 1044 119
rect 559 51 632 67
rect 1086 51 1116 119
rect 1336 66 1366 92
rect 1422 66 1452 92
rect 559 21 1116 51
<< polycont >>
rect 461 426 495 460
rect 103 260 137 294
rect 217 306 251 340
rect 467 318 501 352
rect 359 240 393 274
rect 647 327 681 361
rect 815 327 849 361
rect 926 305 960 339
rect 994 305 1028 339
rect 1211 272 1245 306
rect 582 67 616 101
rect 1211 204 1245 238
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 19 580 89 596
rect 19 546 39 580
rect 73 546 89 580
rect 19 497 89 546
rect 19 463 39 497
rect 73 463 89 497
rect 19 414 89 463
rect 137 580 215 649
rect 137 546 159 580
rect 193 546 215 580
rect 589 580 697 649
rect 137 494 215 546
rect 137 460 159 494
rect 193 460 215 494
rect 137 458 215 460
rect 307 560 481 576
rect 307 526 361 560
rect 395 526 431 560
rect 465 526 481 560
rect 589 546 626 580
rect 660 546 697 580
rect 589 530 697 546
rect 731 580 797 596
rect 731 546 747 580
rect 781 546 797 580
rect 307 510 481 526
rect 307 424 341 510
rect 445 460 511 476
rect 445 444 461 460
rect 19 380 39 414
rect 73 380 89 414
rect 19 364 89 380
rect 123 390 341 424
rect 375 426 461 444
rect 495 444 511 460
rect 731 470 797 546
rect 495 426 665 444
rect 375 410 665 426
rect 19 188 53 364
rect 123 310 157 390
rect 87 294 157 310
rect 87 260 103 294
rect 137 260 157 294
rect 201 340 267 356
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 375 290 409 410
rect 631 377 665 410
rect 731 436 747 470
rect 781 436 797 470
rect 731 420 797 436
rect 842 575 909 591
rect 842 541 859 575
rect 893 541 909 575
rect 842 465 909 541
rect 842 431 859 465
rect 893 431 909 465
rect 87 256 157 260
rect 346 274 409 290
rect 87 222 312 256
rect 346 240 359 274
rect 393 240 409 274
rect 451 352 517 368
rect 451 318 467 352
rect 501 318 517 352
rect 451 277 517 318
rect 631 361 697 377
rect 631 327 647 361
rect 681 327 697 361
rect 631 311 697 327
rect 731 277 765 420
rect 842 415 909 431
rect 943 575 1009 649
rect 943 541 959 575
rect 993 541 1009 575
rect 943 465 1009 541
rect 943 431 959 465
rect 993 431 1009 465
rect 943 415 1009 431
rect 1043 579 1112 591
rect 1043 545 1059 579
rect 1093 545 1112 579
rect 1043 508 1112 545
rect 1043 474 1059 508
rect 1093 474 1112 508
rect 1043 436 1112 474
rect 842 377 876 415
rect 1043 402 1059 436
rect 1093 402 1112 436
rect 1043 390 1112 402
rect 1146 579 1327 649
rect 1146 545 1150 579
rect 1184 545 1277 579
rect 1311 545 1327 579
rect 1146 508 1327 545
rect 1146 474 1150 508
rect 1184 474 1277 508
rect 1311 474 1327 508
rect 1146 440 1327 474
rect 1146 406 1150 440
rect 1184 406 1277 440
rect 1311 406 1327 440
rect 1146 390 1327 406
rect 1361 580 1427 596
rect 1361 546 1373 580
rect 1407 546 1427 580
rect 1361 497 1427 546
rect 1361 463 1373 497
rect 1407 463 1427 497
rect 1361 414 1427 463
rect 799 361 876 377
rect 799 327 815 361
rect 849 327 876 361
rect 799 311 876 327
rect 451 261 807 277
rect 451 243 757 261
rect 346 224 409 240
rect 741 227 757 243
rect 791 227 807 261
rect 278 190 312 222
rect 19 154 244 188
rect 19 146 73 154
rect 19 112 39 146
rect 19 70 73 112
rect 109 86 125 120
rect 159 86 176 120
rect 109 17 176 86
rect 210 85 244 154
rect 278 174 449 190
rect 278 140 380 174
rect 414 140 449 174
rect 584 185 707 201
rect 584 151 600 185
rect 634 151 671 185
rect 705 151 707 185
rect 278 124 449 140
rect 566 101 632 117
rect 566 85 582 101
rect 210 67 582 85
rect 616 67 632 101
rect 210 51 632 67
rect 668 17 707 151
rect 741 171 807 227
rect 741 137 757 171
rect 791 137 807 171
rect 741 121 807 137
rect 842 255 876 311
rect 910 339 1044 356
rect 910 305 926 339
rect 960 305 994 339
rect 1028 305 1044 339
rect 910 289 1044 305
rect 1078 322 1112 390
rect 1361 380 1373 414
rect 1407 380 1427 414
rect 1078 306 1261 322
rect 1078 272 1211 306
rect 1245 272 1261 306
rect 1078 255 1261 272
rect 842 239 919 255
rect 842 205 869 239
rect 903 205 919 239
rect 842 165 919 205
rect 842 131 869 165
rect 903 131 919 165
rect 842 115 919 131
rect 953 239 1019 255
rect 953 205 969 239
rect 1003 205 1019 239
rect 953 165 1019 205
rect 1078 221 1127 255
rect 1161 238 1261 255
rect 1161 221 1211 238
rect 1078 204 1211 221
rect 1245 204 1261 238
rect 1078 188 1261 204
rect 1361 228 1427 380
rect 1463 580 1513 649
rect 1497 546 1513 580
rect 1463 497 1513 546
rect 1497 463 1513 497
rect 1463 414 1513 463
rect 1497 380 1513 414
rect 1463 364 1513 380
rect 1361 194 1377 228
rect 1411 194 1427 228
rect 953 131 969 165
rect 1003 131 1019 165
rect 953 17 1019 131
rect 1111 165 1177 188
rect 1111 131 1127 165
rect 1161 131 1177 165
rect 1111 115 1177 131
rect 1261 138 1327 154
rect 1261 104 1277 138
rect 1311 104 1327 138
rect 1261 17 1327 104
rect 1361 138 1427 194
rect 1361 104 1377 138
rect 1411 104 1427 138
rect 1361 88 1427 104
rect 1463 228 1513 244
rect 1497 194 1513 228
rect 1463 138 1513 194
rect 1497 104 1513 138
rect 1463 17 1513 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel comment s 717 368 717 368 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dlclkp_2
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nbase s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew
flabel corelocali s 1375 94 1409 128 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1375 168 1409 202 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1375 242 1409 276 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1375 390 1409 424 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1375 464 1409 498 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
flabel corelocali s 1375 538 1409 572 0 FreeSans 340 0 0 0 GCLK
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1536 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2909356
string GDS_START 2896962
<< end >>
