magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 101 324 167 370
rect 217 358 317 424
rect 101 290 409 324
rect 359 252 409 290
rect 511 228 553 430
rect 655 236 743 310
rect 2490 364 2541 596
rect 2490 226 2524 364
rect 2425 70 2524 226
rect 2791 70 2858 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 23 492 73 596
rect 113 526 179 649
rect 287 560 389 592
rect 287 526 477 560
rect 511 532 564 649
rect 715 532 781 649
rect 821 581 1162 615
rect 443 498 477 526
rect 821 510 871 581
rect 23 458 409 492
rect 23 256 67 458
rect 359 366 409 458
rect 443 476 759 498
rect 918 476 985 547
rect 443 464 985 476
rect 1024 474 1090 547
rect 23 190 228 256
rect 443 218 477 464
rect 725 442 985 464
rect 587 398 691 430
rect 587 364 843 398
rect 23 70 89 190
rect 301 184 477 218
rect 587 202 621 364
rect 777 244 843 364
rect 123 17 189 156
rect 301 70 367 184
rect 465 17 531 150
rect 587 68 640 202
rect 676 17 742 202
rect 776 85 842 202
rect 884 185 918 442
rect 952 274 1006 408
rect 884 119 938 185
rect 972 85 1006 274
rect 776 51 1006 85
rect 1040 304 1074 474
rect 1128 451 1162 581
rect 1235 485 1285 649
rect 1319 581 1489 615
rect 1319 451 1353 581
rect 1128 417 1353 451
rect 1128 404 1162 417
rect 1108 338 1162 404
rect 1387 383 1421 547
rect 1455 424 1489 581
rect 1523 459 1557 649
rect 1706 581 2076 615
rect 1597 504 1663 551
rect 1706 538 1772 581
rect 1916 504 1966 547
rect 2010 504 2076 581
rect 2116 504 2150 649
rect 2190 504 2256 596
rect 1597 470 1966 504
rect 1597 458 1663 470
rect 1916 458 1966 470
rect 2222 453 2256 504
rect 1809 424 1876 436
rect 2000 424 2256 453
rect 2300 470 2350 596
rect 2390 504 2456 649
rect 2300 436 2447 470
rect 1455 390 1766 424
rect 1210 338 1421 383
rect 1459 350 1525 356
rect 1459 316 1471 350
rect 1505 316 1525 350
rect 1040 270 1422 304
rect 1040 70 1090 270
rect 1345 238 1422 270
rect 1459 249 1525 316
rect 1732 336 1766 390
rect 1809 419 2256 424
rect 1809 390 2034 419
rect 2222 394 2256 419
rect 1809 370 1876 390
rect 1163 181 1297 236
rect 1388 215 1422 238
rect 1567 215 1633 290
rect 1732 270 1798 336
rect 1388 181 1633 215
rect 1842 210 1876 370
rect 2117 356 2183 385
rect 1945 350 2183 356
rect 1945 316 1951 350
rect 1985 316 2183 350
rect 2222 328 2379 394
rect 1945 310 2183 316
rect 2117 251 2183 310
rect 2413 294 2447 436
rect 2245 260 2447 294
rect 1163 147 1354 181
rect 1204 17 1274 113
rect 1320 70 1386 147
rect 1500 17 1659 147
rect 1757 70 1876 210
rect 1924 214 1990 246
rect 2245 214 2279 260
rect 2601 310 2651 575
rect 2691 399 2757 649
rect 2601 244 2757 310
rect 2601 226 2651 244
rect 1924 180 2279 214
rect 2057 17 2179 136
rect 2213 70 2279 180
rect 2325 17 2391 226
rect 2568 108 2651 226
rect 2691 17 2757 210
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 1471 316 1505 350
rect 1951 316 1985 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 1459 350 1517 356
rect 1459 316 1471 350
rect 1505 347 1517 350
rect 1939 350 1997 356
rect 1939 347 1951 350
rect 1505 319 1951 347
rect 1505 316 1517 319
rect 1459 310 1517 316
rect 1939 316 1951 319
rect 1985 316 1997 350
rect 1939 310 1997 316
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
rlabel locali s 217 358 317 424 6 D
port 1 nsew signal input
rlabel locali s 2791 70 2858 596 6 Q
port 2 nsew signal output
rlabel locali s 2490 364 2541 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2490 226 2524 364 6 Q_N
port 3 nsew signal output
rlabel locali s 2425 70 2524 226 6 Q_N
port 3 nsew signal output
rlabel locali s 511 228 553 430 6 SCD
port 4 nsew signal input
rlabel locali s 359 252 409 290 6 SCE
port 5 nsew signal input
rlabel locali s 101 324 167 370 6 SCE
port 5 nsew signal input
rlabel locali s 101 290 409 324 6 SCE
port 5 nsew signal input
rlabel metal1 s 1939 347 1997 356 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1939 310 1997 319 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1459 347 1517 356 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1459 319 1997 347 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1459 310 1517 319 6 SET_B
port 6 nsew signal input
rlabel locali s 655 236 743 310 6 CLK
port 7 nsew clock input
rlabel metal1 s 0 -49 2880 49 8 VGND
port 8 nsew ground bidirectional
rlabel metal1 s 0 617 2880 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 172610
string GDS_START 151162
<< end >>
