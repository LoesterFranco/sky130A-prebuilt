magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 93 47 123 177
rect 187 47 217 177
rect 271 47 301 177
rect 453 47 483 177
rect 557 47 587 177
rect 681 47 711 177
rect 765 47 795 177
rect 883 47 913 177
<< pmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 579 297 615 497
rect 673 297 709 497
rect 767 297 803 497
rect 885 297 921 497
<< ndiff >>
rect 27 157 93 177
rect 27 123 39 157
rect 73 123 93 157
rect 27 89 93 123
rect 27 55 39 89
rect 73 55 93 89
rect 27 47 93 55
rect 123 93 187 177
rect 123 59 133 93
rect 167 59 187 93
rect 123 47 187 59
rect 217 157 271 177
rect 217 123 227 157
rect 261 123 271 157
rect 217 89 271 123
rect 217 55 227 89
rect 261 55 271 89
rect 217 47 271 55
rect 301 93 453 177
rect 301 59 321 93
rect 355 59 389 93
rect 423 59 453 93
rect 301 47 453 59
rect 483 157 557 177
rect 483 123 501 157
rect 535 123 557 157
rect 483 89 557 123
rect 483 55 501 89
rect 535 55 557 89
rect 483 47 557 55
rect 587 89 681 177
rect 587 55 611 89
rect 645 55 681 89
rect 587 47 681 55
rect 711 157 765 177
rect 711 123 721 157
rect 755 123 765 157
rect 711 89 765 123
rect 711 55 721 89
rect 755 55 765 89
rect 711 47 765 55
rect 795 168 883 177
rect 795 134 831 168
rect 865 134 883 168
rect 795 47 883 134
rect 913 101 976 177
rect 913 67 934 101
rect 968 67 976 101
rect 913 47 976 67
<< pdiff >>
rect 27 489 85 497
rect 27 455 39 489
rect 73 455 85 489
rect 27 421 85 455
rect 27 387 39 421
rect 73 387 85 421
rect 27 353 85 387
rect 27 319 39 353
rect 73 319 85 353
rect 27 297 85 319
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 417 179 451
rect 121 383 133 417
rect 167 383 179 417
rect 121 297 179 383
rect 215 489 273 497
rect 215 455 227 489
rect 261 455 273 489
rect 215 421 273 455
rect 215 387 227 421
rect 261 387 273 421
rect 215 353 273 387
rect 215 319 227 353
rect 261 319 273 353
rect 215 297 273 319
rect 309 444 367 497
rect 309 410 321 444
rect 355 410 367 444
rect 309 297 367 410
rect 403 421 457 497
rect 403 387 415 421
rect 449 387 457 421
rect 403 353 457 387
rect 403 319 415 353
rect 449 319 457 353
rect 403 297 457 319
rect 521 421 579 497
rect 521 387 533 421
rect 567 387 579 421
rect 521 353 579 387
rect 521 319 533 353
rect 567 319 579 353
rect 521 297 579 319
rect 615 444 673 497
rect 615 410 627 444
rect 661 410 673 444
rect 615 297 673 410
rect 709 489 767 497
rect 709 455 721 489
rect 755 455 767 489
rect 709 421 767 455
rect 709 387 721 421
rect 755 387 767 421
rect 709 353 767 387
rect 709 319 721 353
rect 755 319 767 353
rect 709 297 767 319
rect 803 489 885 497
rect 803 455 831 489
rect 865 455 885 489
rect 803 421 885 455
rect 803 387 831 421
rect 865 387 885 421
rect 803 297 885 387
rect 921 438 975 497
rect 921 404 933 438
rect 967 404 975 438
rect 921 370 975 404
rect 921 336 933 370
rect 967 336 975 370
rect 921 297 975 336
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 133 59 167 93
rect 227 123 261 157
rect 227 55 261 89
rect 321 59 355 93
rect 389 59 423 93
rect 501 123 535 157
rect 501 55 535 89
rect 611 55 645 89
rect 721 123 755 157
rect 721 55 755 89
rect 831 134 865 168
rect 934 67 968 101
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 39 319 73 353
rect 133 451 167 485
rect 133 383 167 417
rect 227 455 261 489
rect 227 387 261 421
rect 227 319 261 353
rect 321 410 355 444
rect 415 387 449 421
rect 415 319 449 353
rect 533 387 567 421
rect 533 319 567 353
rect 627 410 661 444
rect 721 455 755 489
rect 721 387 755 421
rect 721 319 755 353
rect 831 455 865 489
rect 831 387 865 421
rect 933 404 967 438
rect 933 336 967 370
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 579 497 615 523
rect 673 497 709 523
rect 767 497 803 523
rect 885 497 921 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 579 282 615 297
rect 673 282 709 297
rect 767 282 803 297
rect 885 282 921 297
rect 83 259 123 282
rect 177 259 217 282
rect 63 249 217 259
rect 63 215 79 249
rect 113 215 157 249
rect 191 215 217 249
rect 63 205 217 215
rect 93 177 123 205
rect 187 177 217 205
rect 271 259 311 282
rect 365 259 405 282
rect 577 259 617 282
rect 671 259 711 282
rect 271 249 483 259
rect 271 215 328 249
rect 362 215 406 249
rect 440 215 483 249
rect 271 205 483 215
rect 271 177 301 205
rect 453 177 483 205
rect 557 249 711 259
rect 557 215 573 249
rect 607 215 651 249
rect 685 215 711 249
rect 557 205 711 215
rect 557 177 587 205
rect 681 177 711 205
rect 765 265 805 282
rect 883 265 923 282
rect 765 249 989 265
rect 765 215 945 249
rect 979 215 989 249
rect 765 199 989 215
rect 765 177 795 199
rect 883 177 913 199
rect 93 21 123 47
rect 187 21 217 47
rect 271 21 301 47
rect 453 21 483 47
rect 557 21 587 47
rect 681 21 711 47
rect 765 21 795 47
rect 883 21 913 47
<< polycont >>
rect 79 215 113 249
rect 157 215 191 249
rect 328 215 362 249
rect 406 215 440 249
rect 573 215 607 249
rect 651 215 685 249
rect 945 215 979 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 18 489 89 493
rect 18 455 39 489
rect 73 455 89 489
rect 18 421 89 455
rect 18 387 39 421
rect 73 387 89 421
rect 18 353 89 387
rect 133 485 167 527
rect 133 417 167 451
rect 133 367 167 383
rect 201 489 277 493
rect 201 455 227 489
rect 261 455 277 489
rect 201 421 277 455
rect 201 387 227 421
rect 261 387 277 421
rect 18 319 39 353
rect 73 333 89 353
rect 201 353 277 387
rect 321 459 661 493
rect 321 444 355 459
rect 627 444 661 459
rect 321 367 355 410
rect 389 421 465 425
rect 389 387 415 421
rect 449 387 465 421
rect 201 333 227 353
rect 73 319 227 333
rect 261 333 277 353
rect 389 353 465 387
rect 389 333 415 353
rect 261 319 415 333
rect 449 319 465 353
rect 18 299 465 319
rect 517 421 583 425
rect 517 387 533 421
rect 567 387 583 421
rect 517 353 583 387
rect 627 367 661 410
rect 695 489 771 493
rect 695 455 721 489
rect 755 455 771 489
rect 695 421 771 455
rect 695 387 721 421
rect 755 387 771 421
rect 517 319 533 353
rect 567 333 583 353
rect 695 353 771 387
rect 815 489 881 527
rect 815 455 831 489
rect 865 455 881 489
rect 815 421 881 455
rect 815 387 831 421
rect 865 387 881 421
rect 815 367 881 387
rect 925 438 993 493
rect 925 404 933 438
rect 967 404 993 438
rect 925 370 993 404
rect 695 333 721 353
rect 567 319 721 333
rect 755 333 771 353
rect 925 336 933 370
rect 967 336 993 370
rect 925 333 993 336
rect 755 319 993 333
rect 517 299 993 319
rect 18 249 262 265
rect 18 215 79 249
rect 113 215 157 249
rect 191 215 262 249
rect 18 211 262 215
rect 300 249 484 265
rect 300 215 328 249
rect 362 215 406 249
rect 440 215 484 249
rect 300 211 484 215
rect 540 249 711 265
rect 540 215 573 249
rect 607 215 651 249
rect 685 215 711 249
rect 540 211 711 215
rect 18 157 771 177
rect 18 123 39 157
rect 73 143 227 157
rect 73 123 89 143
rect 18 89 89 123
rect 201 123 227 143
rect 261 143 501 157
rect 261 123 277 143
rect 18 55 39 89
rect 73 55 89 89
rect 18 51 89 55
rect 133 93 167 109
rect 133 17 167 59
rect 201 89 277 123
rect 485 123 501 143
rect 535 143 721 157
rect 535 123 551 143
rect 201 55 227 89
rect 261 55 277 89
rect 201 51 277 55
rect 321 93 433 109
rect 355 59 389 93
rect 423 59 433 93
rect 321 17 433 59
rect 485 89 551 123
rect 695 123 721 143
rect 755 123 771 157
rect 485 55 501 89
rect 535 55 551 89
rect 485 51 551 55
rect 585 89 661 109
rect 585 55 611 89
rect 645 55 661 89
rect 585 17 661 55
rect 695 89 771 123
rect 815 168 891 299
rect 815 134 831 168
rect 865 134 891 168
rect 926 249 994 265
rect 926 215 945 249
rect 979 215 994 249
rect 926 151 994 215
rect 815 119 891 134
rect 695 55 721 89
rect 755 85 771 89
rect 926 101 993 117
rect 926 85 934 101
rect 755 67 934 85
rect 968 67 993 101
rect 755 55 993 67
rect 695 51 993 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel corelocali s 132 221 166 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel corelocali s 948 425 982 459 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 846 289 880 323 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 846 221 880 255 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 540 357 574 391 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 948 357 982 391 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 846 153 880 187 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel corelocali s 948 153 982 187 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 947 221 981 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel corelocali s 671 221 705 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 580 221 614 255 0 FreeSans 200 0 0 0 A3
port 3 nsew
flabel corelocali s 397 221 431 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 310 221 344 255 0 FreeSans 200 0 0 0 A2
port 2 nsew
flabel corelocali s 215 221 249 255 0 FreeSans 200 0 0 0 A1
port 1 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 o31ai_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 559036
string GDS_START 549708
<< end >>
