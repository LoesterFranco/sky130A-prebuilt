magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 332 2438 704
<< pwell >>
rect 0 0 2400 49
<< scnmos >>
rect 84 74 114 222
rect 182 74 212 222
rect 268 74 298 222
rect 354 74 384 222
rect 440 74 470 222
rect 526 74 556 222
rect 612 74 642 222
rect 712 74 742 222
rect 798 74 828 222
rect 898 74 928 222
rect 984 74 1014 222
rect 1070 74 1100 222
rect 1156 74 1186 222
rect 1256 74 1286 222
rect 1342 74 1372 222
rect 1442 74 1472 222
rect 1528 74 1558 222
rect 1628 74 1658 222
rect 1714 74 1744 222
rect 1814 74 1844 222
rect 1900 74 1930 222
rect 2000 74 2030 222
rect 2086 74 2116 222
rect 2186 74 2216 222
rect 2272 74 2302 222
<< pmoshvt >>
rect 87 368 117 592
rect 177 368 207 592
rect 267 368 297 592
rect 357 368 387 592
rect 451 368 481 592
rect 541 368 571 592
rect 631 368 661 592
rect 721 368 751 592
rect 811 368 841 592
rect 901 368 931 592
rect 991 368 1021 592
rect 1081 368 1111 592
rect 1171 368 1201 592
rect 1261 368 1291 592
rect 1351 368 1381 592
rect 1441 368 1471 592
rect 1531 368 1561 592
rect 1621 368 1651 592
rect 1711 368 1741 592
rect 1811 368 1841 592
rect 1901 368 1931 592
rect 2001 368 2031 592
rect 2091 368 2121 592
rect 2183 368 2213 592
rect 2281 368 2311 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 152 182 222
rect 114 118 125 152
rect 159 118 182 152
rect 114 74 182 118
rect 212 210 268 222
rect 212 176 223 210
rect 257 176 268 210
rect 212 120 268 176
rect 212 86 223 120
rect 257 86 268 120
rect 212 74 268 86
rect 298 152 354 222
rect 298 118 309 152
rect 343 118 354 152
rect 298 74 354 118
rect 384 210 440 222
rect 384 176 395 210
rect 429 176 440 210
rect 384 120 440 176
rect 384 86 395 120
rect 429 86 440 120
rect 384 74 440 86
rect 470 142 526 222
rect 470 108 481 142
rect 515 108 526 142
rect 470 74 526 108
rect 556 210 612 222
rect 556 176 567 210
rect 601 176 612 210
rect 556 120 612 176
rect 556 86 567 120
rect 601 86 612 120
rect 556 74 612 86
rect 642 142 712 222
rect 642 108 653 142
rect 687 108 712 142
rect 642 74 712 108
rect 742 210 798 222
rect 742 176 753 210
rect 787 176 798 210
rect 742 120 798 176
rect 742 86 753 120
rect 787 86 798 120
rect 742 74 798 86
rect 828 210 898 222
rect 828 176 839 210
rect 873 176 898 210
rect 828 120 898 176
rect 828 86 839 120
rect 873 86 898 120
rect 828 74 898 86
rect 928 210 984 222
rect 928 176 939 210
rect 973 176 984 210
rect 928 120 984 176
rect 928 86 939 120
rect 973 86 984 120
rect 928 74 984 86
rect 1014 205 1070 222
rect 1014 171 1025 205
rect 1059 171 1070 205
rect 1014 120 1070 171
rect 1014 86 1025 120
rect 1059 86 1070 120
rect 1014 74 1070 86
rect 1100 210 1156 222
rect 1100 176 1111 210
rect 1145 176 1156 210
rect 1100 120 1156 176
rect 1100 86 1111 120
rect 1145 86 1156 120
rect 1100 74 1156 86
rect 1186 205 1256 222
rect 1186 171 1197 205
rect 1231 171 1256 205
rect 1186 120 1256 171
rect 1186 86 1197 120
rect 1231 86 1256 120
rect 1186 74 1256 86
rect 1286 210 1342 222
rect 1286 176 1297 210
rect 1331 176 1342 210
rect 1286 120 1342 176
rect 1286 86 1297 120
rect 1331 86 1342 120
rect 1286 74 1342 86
rect 1372 205 1442 222
rect 1372 171 1383 205
rect 1417 171 1442 205
rect 1372 120 1442 171
rect 1372 86 1383 120
rect 1417 86 1442 120
rect 1372 74 1442 86
rect 1472 210 1528 222
rect 1472 176 1483 210
rect 1517 176 1528 210
rect 1472 120 1528 176
rect 1472 86 1483 120
rect 1517 86 1528 120
rect 1472 74 1528 86
rect 1558 205 1628 222
rect 1558 171 1569 205
rect 1603 171 1628 205
rect 1558 120 1628 171
rect 1558 86 1569 120
rect 1603 86 1628 120
rect 1558 74 1628 86
rect 1658 210 1714 222
rect 1658 176 1669 210
rect 1703 176 1714 210
rect 1658 120 1714 176
rect 1658 86 1669 120
rect 1703 86 1714 120
rect 1658 74 1714 86
rect 1744 205 1814 222
rect 1744 171 1755 205
rect 1789 171 1814 205
rect 1744 120 1814 171
rect 1744 86 1755 120
rect 1789 86 1814 120
rect 1744 74 1814 86
rect 1844 210 1900 222
rect 1844 176 1855 210
rect 1889 176 1900 210
rect 1844 120 1900 176
rect 1844 86 1855 120
rect 1889 86 1900 120
rect 1844 74 1900 86
rect 1930 205 2000 222
rect 1930 171 1941 205
rect 1975 171 2000 205
rect 1930 120 2000 171
rect 1930 86 1941 120
rect 1975 86 2000 120
rect 1930 74 2000 86
rect 2030 210 2086 222
rect 2030 176 2041 210
rect 2075 176 2086 210
rect 2030 120 2086 176
rect 2030 86 2041 120
rect 2075 86 2086 120
rect 2030 74 2086 86
rect 2116 205 2186 222
rect 2116 171 2127 205
rect 2161 171 2186 205
rect 2116 120 2186 171
rect 2116 86 2127 120
rect 2161 86 2186 120
rect 2116 74 2186 86
rect 2216 210 2272 222
rect 2216 176 2227 210
rect 2261 176 2272 210
rect 2216 120 2272 176
rect 2216 86 2227 120
rect 2261 86 2272 120
rect 2216 74 2272 86
rect 2302 210 2373 222
rect 2302 176 2327 210
rect 2361 176 2373 210
rect 2302 120 2373 176
rect 2302 86 2327 120
rect 2361 86 2373 120
rect 2302 74 2373 86
<< pdiff >>
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 510 87 546
rect 28 476 40 510
rect 74 476 87 510
rect 28 440 87 476
rect 28 406 40 440
rect 74 406 87 440
rect 28 368 87 406
rect 117 580 177 592
rect 117 546 130 580
rect 164 546 177 580
rect 117 508 177 546
rect 117 474 130 508
rect 164 474 177 508
rect 117 368 177 474
rect 207 580 267 592
rect 207 546 220 580
rect 254 546 267 580
rect 207 510 267 546
rect 207 476 220 510
rect 254 476 267 510
rect 207 440 267 476
rect 207 406 220 440
rect 254 406 267 440
rect 207 368 267 406
rect 297 580 357 592
rect 297 546 310 580
rect 344 546 357 580
rect 297 508 357 546
rect 297 474 310 508
rect 344 474 357 508
rect 297 368 357 474
rect 387 580 451 592
rect 387 546 404 580
rect 438 546 451 580
rect 387 497 451 546
rect 387 463 404 497
rect 438 463 451 497
rect 387 414 451 463
rect 387 380 404 414
rect 438 380 451 414
rect 387 368 451 380
rect 481 580 541 592
rect 481 546 494 580
rect 528 546 541 580
rect 481 478 541 546
rect 481 444 494 478
rect 528 444 541 478
rect 481 368 541 444
rect 571 580 631 592
rect 571 546 584 580
rect 618 546 631 580
rect 571 497 631 546
rect 571 463 584 497
rect 618 463 631 497
rect 571 414 631 463
rect 571 380 584 414
rect 618 380 631 414
rect 571 368 631 380
rect 661 580 721 592
rect 661 546 674 580
rect 708 546 721 580
rect 661 478 721 546
rect 661 444 674 478
rect 708 444 721 478
rect 661 368 721 444
rect 751 580 811 592
rect 751 546 764 580
rect 798 546 811 580
rect 751 497 811 546
rect 751 463 764 497
rect 798 463 811 497
rect 751 414 811 463
rect 751 380 764 414
rect 798 380 811 414
rect 751 368 811 380
rect 841 580 901 592
rect 841 546 854 580
rect 888 546 901 580
rect 841 506 901 546
rect 841 472 854 506
rect 888 472 901 506
rect 841 434 901 472
rect 841 400 854 434
rect 888 400 901 434
rect 841 368 901 400
rect 931 580 991 592
rect 931 546 944 580
rect 978 546 991 580
rect 931 497 991 546
rect 931 463 944 497
rect 978 463 991 497
rect 931 418 991 463
rect 931 384 944 418
rect 978 384 991 418
rect 931 368 991 384
rect 1021 580 1081 592
rect 1021 546 1034 580
rect 1068 546 1081 580
rect 1021 506 1081 546
rect 1021 472 1034 506
rect 1068 472 1081 506
rect 1021 434 1081 472
rect 1021 400 1034 434
rect 1068 400 1081 434
rect 1021 368 1081 400
rect 1111 580 1171 592
rect 1111 546 1124 580
rect 1158 546 1171 580
rect 1111 497 1171 546
rect 1111 463 1124 497
rect 1158 463 1171 497
rect 1111 418 1171 463
rect 1111 384 1124 418
rect 1158 384 1171 418
rect 1111 368 1171 384
rect 1201 580 1261 592
rect 1201 546 1214 580
rect 1248 546 1261 580
rect 1201 506 1261 546
rect 1201 472 1214 506
rect 1248 472 1261 506
rect 1201 434 1261 472
rect 1201 400 1214 434
rect 1248 400 1261 434
rect 1201 368 1261 400
rect 1291 580 1351 592
rect 1291 546 1304 580
rect 1338 546 1351 580
rect 1291 497 1351 546
rect 1291 463 1304 497
rect 1338 463 1351 497
rect 1291 418 1351 463
rect 1291 384 1304 418
rect 1338 384 1351 418
rect 1291 368 1351 384
rect 1381 580 1441 592
rect 1381 546 1394 580
rect 1428 546 1441 580
rect 1381 506 1441 546
rect 1381 472 1394 506
rect 1428 472 1441 506
rect 1381 434 1441 472
rect 1381 400 1394 434
rect 1428 400 1441 434
rect 1381 368 1441 400
rect 1471 580 1531 592
rect 1471 546 1484 580
rect 1518 546 1531 580
rect 1471 497 1531 546
rect 1471 463 1484 497
rect 1518 463 1531 497
rect 1471 418 1531 463
rect 1471 384 1484 418
rect 1518 384 1531 418
rect 1471 368 1531 384
rect 1561 580 1621 592
rect 1561 546 1574 580
rect 1608 546 1621 580
rect 1561 506 1621 546
rect 1561 472 1574 506
rect 1608 472 1621 506
rect 1561 434 1621 472
rect 1561 400 1574 434
rect 1608 400 1621 434
rect 1561 368 1621 400
rect 1651 580 1711 592
rect 1651 546 1664 580
rect 1698 546 1711 580
rect 1651 497 1711 546
rect 1651 463 1664 497
rect 1698 463 1711 497
rect 1651 414 1711 463
rect 1651 380 1664 414
rect 1698 380 1711 414
rect 1651 368 1711 380
rect 1741 580 1811 592
rect 1741 546 1754 580
rect 1788 546 1811 580
rect 1741 506 1811 546
rect 1741 472 1754 506
rect 1788 472 1811 506
rect 1741 434 1811 472
rect 1741 400 1754 434
rect 1788 400 1811 434
rect 1741 368 1811 400
rect 1841 580 1901 592
rect 1841 546 1854 580
rect 1888 546 1901 580
rect 1841 497 1901 546
rect 1841 463 1854 497
rect 1888 463 1901 497
rect 1841 414 1901 463
rect 1841 380 1854 414
rect 1888 380 1901 414
rect 1841 368 1901 380
rect 1931 580 2001 592
rect 1931 546 1944 580
rect 1978 546 2001 580
rect 1931 506 2001 546
rect 1931 472 1944 506
rect 1978 472 2001 506
rect 1931 434 2001 472
rect 1931 400 1944 434
rect 1978 400 2001 434
rect 1931 368 2001 400
rect 2031 580 2091 592
rect 2031 546 2044 580
rect 2078 546 2091 580
rect 2031 497 2091 546
rect 2031 463 2044 497
rect 2078 463 2091 497
rect 2031 418 2091 463
rect 2031 384 2044 418
rect 2078 384 2091 418
rect 2031 368 2091 384
rect 2121 580 2183 592
rect 2121 546 2134 580
rect 2168 546 2183 580
rect 2121 506 2183 546
rect 2121 472 2134 506
rect 2168 472 2183 506
rect 2121 434 2183 472
rect 2121 400 2134 434
rect 2168 400 2183 434
rect 2121 368 2183 400
rect 2213 580 2281 592
rect 2213 546 2234 580
rect 2268 546 2281 580
rect 2213 497 2281 546
rect 2213 463 2234 497
rect 2268 463 2281 497
rect 2213 414 2281 463
rect 2213 380 2234 414
rect 2268 380 2281 414
rect 2213 368 2281 380
rect 2311 580 2370 592
rect 2311 546 2324 580
rect 2358 546 2370 580
rect 2311 497 2370 546
rect 2311 463 2324 497
rect 2358 463 2370 497
rect 2311 414 2370 463
rect 2311 380 2324 414
rect 2358 380 2370 414
rect 2311 368 2370 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 118 159 152
rect 223 176 257 210
rect 223 86 257 120
rect 309 118 343 152
rect 395 176 429 210
rect 395 86 429 120
rect 481 108 515 142
rect 567 176 601 210
rect 567 86 601 120
rect 653 108 687 142
rect 753 176 787 210
rect 753 86 787 120
rect 839 176 873 210
rect 839 86 873 120
rect 939 176 973 210
rect 939 86 973 120
rect 1025 171 1059 205
rect 1025 86 1059 120
rect 1111 176 1145 210
rect 1111 86 1145 120
rect 1197 171 1231 205
rect 1197 86 1231 120
rect 1297 176 1331 210
rect 1297 86 1331 120
rect 1383 171 1417 205
rect 1383 86 1417 120
rect 1483 176 1517 210
rect 1483 86 1517 120
rect 1569 171 1603 205
rect 1569 86 1603 120
rect 1669 176 1703 210
rect 1669 86 1703 120
rect 1755 171 1789 205
rect 1755 86 1789 120
rect 1855 176 1889 210
rect 1855 86 1889 120
rect 1941 171 1975 205
rect 1941 86 1975 120
rect 2041 176 2075 210
rect 2041 86 2075 120
rect 2127 171 2161 205
rect 2127 86 2161 120
rect 2227 176 2261 210
rect 2227 86 2261 120
rect 2327 176 2361 210
rect 2327 86 2361 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 474 164 508
rect 220 546 254 580
rect 220 476 254 510
rect 220 406 254 440
rect 310 546 344 580
rect 310 474 344 508
rect 404 546 438 580
rect 404 463 438 497
rect 404 380 438 414
rect 494 546 528 580
rect 494 444 528 478
rect 584 546 618 580
rect 584 463 618 497
rect 584 380 618 414
rect 674 546 708 580
rect 674 444 708 478
rect 764 546 798 580
rect 764 463 798 497
rect 764 380 798 414
rect 854 546 888 580
rect 854 472 888 506
rect 854 400 888 434
rect 944 546 978 580
rect 944 463 978 497
rect 944 384 978 418
rect 1034 546 1068 580
rect 1034 472 1068 506
rect 1034 400 1068 434
rect 1124 546 1158 580
rect 1124 463 1158 497
rect 1124 384 1158 418
rect 1214 546 1248 580
rect 1214 472 1248 506
rect 1214 400 1248 434
rect 1304 546 1338 580
rect 1304 463 1338 497
rect 1304 384 1338 418
rect 1394 546 1428 580
rect 1394 472 1428 506
rect 1394 400 1428 434
rect 1484 546 1518 580
rect 1484 463 1518 497
rect 1484 384 1518 418
rect 1574 546 1608 580
rect 1574 472 1608 506
rect 1574 400 1608 434
rect 1664 546 1698 580
rect 1664 463 1698 497
rect 1664 380 1698 414
rect 1754 546 1788 580
rect 1754 472 1788 506
rect 1754 400 1788 434
rect 1854 546 1888 580
rect 1854 463 1888 497
rect 1854 380 1888 414
rect 1944 546 1978 580
rect 1944 472 1978 506
rect 1944 400 1978 434
rect 2044 546 2078 580
rect 2044 463 2078 497
rect 2044 384 2078 418
rect 2134 546 2168 580
rect 2134 472 2168 506
rect 2134 400 2168 434
rect 2234 546 2268 580
rect 2234 463 2268 497
rect 2234 380 2268 414
rect 2324 546 2358 580
rect 2324 463 2358 497
rect 2324 380 2358 414
<< poly >>
rect 87 592 117 618
rect 177 592 207 618
rect 267 592 297 618
rect 357 592 387 618
rect 451 592 481 618
rect 541 592 571 618
rect 631 592 661 618
rect 721 592 751 618
rect 811 592 841 618
rect 901 592 931 618
rect 991 592 1021 618
rect 1081 592 1111 618
rect 1171 592 1201 618
rect 1261 592 1291 618
rect 1351 592 1381 618
rect 1441 592 1471 618
rect 1531 592 1561 618
rect 1621 592 1651 618
rect 1711 592 1741 618
rect 1811 592 1841 618
rect 1901 592 1931 618
rect 2001 592 2031 618
rect 2091 592 2121 618
rect 2183 592 2213 618
rect 2281 592 2311 618
rect 87 353 117 368
rect 177 353 207 368
rect 267 353 297 368
rect 357 353 387 368
rect 451 353 481 368
rect 541 353 571 368
rect 631 353 661 368
rect 721 353 751 368
rect 811 353 841 368
rect 901 353 931 368
rect 991 353 1021 368
rect 1081 353 1111 368
rect 1171 353 1201 368
rect 1261 353 1291 368
rect 1351 353 1381 368
rect 1441 353 1471 368
rect 1531 353 1561 368
rect 1621 353 1651 368
rect 1711 353 1741 368
rect 1811 353 1841 368
rect 1901 353 1931 368
rect 2001 353 2031 368
rect 2091 353 2121 368
rect 2183 353 2213 368
rect 2281 353 2311 368
rect 84 336 120 353
rect 174 336 210 353
rect 264 336 300 353
rect 84 320 300 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 300 320
rect 84 270 300 286
rect 354 326 390 353
rect 448 326 484 353
rect 538 326 574 353
rect 628 326 664 353
rect 718 326 754 353
rect 354 310 754 326
rect 354 276 370 310
rect 404 276 438 310
rect 472 276 506 310
rect 540 276 574 310
rect 608 276 642 310
rect 676 290 754 310
rect 808 290 844 353
rect 676 276 844 290
rect 84 222 114 270
rect 182 222 212 270
rect 268 222 298 270
rect 354 260 844 276
rect 898 326 934 353
rect 988 326 1024 353
rect 1078 326 1114 353
rect 1168 326 1204 353
rect 1258 326 1294 353
rect 1348 326 1384 353
rect 1438 326 1474 353
rect 1528 326 1564 353
rect 1618 326 1654 353
rect 1708 326 1744 353
rect 1808 326 1844 353
rect 1898 326 1934 353
rect 1998 326 2034 353
rect 2088 326 2124 353
rect 2180 326 2216 353
rect 2278 326 2314 353
rect 898 310 2314 326
rect 898 276 1018 310
rect 1052 276 1196 310
rect 1230 276 1384 310
rect 1418 276 1568 310
rect 1602 276 1753 310
rect 1787 276 1939 310
rect 1973 276 2125 310
rect 2159 276 2314 310
rect 898 260 2314 276
rect 354 222 384 260
rect 440 222 470 260
rect 526 222 556 260
rect 612 222 642 260
rect 712 222 742 260
rect 798 222 828 260
rect 898 222 928 260
rect 984 222 1014 260
rect 1070 222 1100 260
rect 1156 222 1186 260
rect 1256 222 1286 260
rect 1342 222 1372 260
rect 1442 222 1472 260
rect 1528 222 1558 260
rect 1628 222 1658 260
rect 1714 222 1744 260
rect 1814 222 1844 260
rect 1900 222 1930 260
rect 2000 222 2030 260
rect 2086 222 2116 260
rect 2186 222 2216 260
rect 2272 222 2302 260
rect 84 48 114 74
rect 182 48 212 74
rect 268 48 298 74
rect 354 48 384 74
rect 440 48 470 74
rect 526 48 556 74
rect 612 48 642 74
rect 712 48 742 74
rect 798 48 828 74
rect 898 48 928 74
rect 984 48 1014 74
rect 1070 48 1100 74
rect 1156 48 1186 74
rect 1256 48 1286 74
rect 1342 48 1372 74
rect 1442 48 1472 74
rect 1528 48 1558 74
rect 1628 48 1658 74
rect 1714 48 1744 74
rect 1814 48 1844 74
rect 1900 48 1930 74
rect 2000 48 2030 74
rect 2086 48 2116 74
rect 2186 48 2216 74
rect 2272 48 2302 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 370 276 404 310
rect 438 276 472 310
rect 506 276 540 310
rect 574 276 608 310
rect 642 276 676 310
rect 1018 276 1052 310
rect 1196 276 1230 310
rect 1384 276 1418 310
rect 1568 276 1602 310
rect 1753 276 1787 310
rect 1939 276 1973 310
rect 2125 276 2159 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 24 580 90 596
rect 24 546 40 580
rect 74 546 90 580
rect 24 510 90 546
rect 24 476 40 510
rect 74 476 90 510
rect 24 440 90 476
rect 130 580 164 649
rect 130 508 164 546
rect 130 458 164 474
rect 204 580 270 596
rect 204 546 220 580
rect 254 546 270 580
rect 204 510 270 546
rect 204 476 220 510
rect 254 476 270 510
rect 24 406 40 440
rect 74 424 90 440
rect 204 440 270 476
rect 310 580 344 649
rect 310 508 344 546
rect 310 458 344 474
rect 388 580 454 596
rect 388 546 404 580
rect 438 546 454 580
rect 388 497 454 546
rect 388 463 404 497
rect 438 463 454 497
rect 204 424 220 440
rect 74 406 220 424
rect 254 424 270 440
rect 254 406 354 424
rect 24 390 354 406
rect 25 320 286 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 286 320
rect 25 270 286 286
rect 320 326 354 390
rect 388 414 454 463
rect 494 580 528 649
rect 494 478 528 546
rect 494 428 528 444
rect 568 580 634 596
rect 568 546 584 580
rect 618 546 634 580
rect 568 497 634 546
rect 568 463 584 497
rect 618 463 634 497
rect 388 380 404 414
rect 438 394 454 414
rect 568 414 634 463
rect 674 580 708 649
rect 674 478 708 546
rect 674 428 708 444
rect 748 580 814 596
rect 748 546 764 580
rect 798 546 814 580
rect 748 497 814 546
rect 748 463 764 497
rect 798 463 814 497
rect 568 394 584 414
rect 438 380 584 394
rect 618 394 634 414
rect 748 414 814 463
rect 748 394 764 414
rect 618 380 764 394
rect 798 380 814 414
rect 854 580 888 649
rect 854 506 888 546
rect 854 434 888 472
rect 928 580 994 596
rect 928 546 944 580
rect 978 546 994 580
rect 928 497 994 546
rect 928 463 944 497
rect 978 463 994 497
rect 928 424 994 463
rect 928 418 946 424
rect 928 404 944 418
rect 854 384 888 400
rect 923 384 944 404
rect 980 390 994 424
rect 978 384 994 390
rect 1034 580 1068 649
rect 1034 506 1068 546
rect 1034 434 1068 472
rect 1108 580 1174 596
rect 1108 546 1124 580
rect 1158 546 1174 580
rect 1108 497 1174 546
rect 1108 463 1124 497
rect 1158 463 1174 497
rect 1108 424 1174 463
rect 1108 404 1124 424
rect 1034 384 1068 400
rect 1102 384 1124 404
rect 1158 384 1174 424
rect 1214 580 1248 649
rect 1214 506 1248 546
rect 1214 434 1248 472
rect 1288 580 1354 596
rect 1288 546 1304 580
rect 1338 546 1354 580
rect 1288 497 1354 546
rect 1288 463 1304 497
rect 1338 463 1354 497
rect 1288 424 1354 463
rect 1288 404 1304 424
rect 1214 384 1248 400
rect 1284 384 1304 404
rect 1338 384 1354 424
rect 1394 580 1428 649
rect 1394 506 1428 546
rect 1394 434 1428 472
rect 1394 384 1428 400
rect 1468 580 1534 596
rect 1468 546 1484 580
rect 1518 546 1534 580
rect 1468 497 1534 546
rect 1468 463 1484 497
rect 1518 463 1534 497
rect 1468 424 1534 463
rect 1468 384 1484 424
rect 1518 384 1534 424
rect 1574 580 1608 649
rect 1574 506 1608 546
rect 1574 434 1608 472
rect 1648 580 1714 596
rect 1648 546 1664 580
rect 1698 546 1714 580
rect 1648 497 1714 546
rect 1648 463 1664 497
rect 1698 463 1714 497
rect 1648 424 1714 463
rect 1648 404 1664 424
rect 1574 384 1608 400
rect 388 360 814 380
rect 748 350 814 360
rect 320 310 692 326
rect 320 276 370 310
rect 404 276 438 310
rect 472 276 506 310
rect 540 276 574 310
rect 608 276 642 310
rect 676 276 692 310
rect 320 260 692 276
rect 748 316 845 350
rect 879 316 887 350
rect 748 260 887 316
rect 320 236 354 260
rect 23 210 354 236
rect 737 226 787 260
rect 23 176 39 210
rect 73 202 223 210
rect 23 120 73 176
rect 257 202 354 210
rect 395 210 787 226
rect 23 86 39 120
rect 23 70 73 86
rect 109 152 175 168
rect 109 118 125 152
rect 159 118 175 152
rect 109 17 175 118
rect 223 120 257 176
rect 429 192 567 210
rect 223 70 257 86
rect 293 152 359 168
rect 293 118 309 152
rect 343 118 359 152
rect 293 17 359 118
rect 395 120 429 176
rect 551 176 567 192
rect 601 192 753 210
rect 395 70 429 86
rect 465 142 515 158
rect 465 108 481 142
rect 465 17 515 108
rect 551 120 601 176
rect 737 176 753 192
rect 551 86 567 120
rect 551 70 601 86
rect 637 142 703 158
rect 637 108 653 142
rect 687 108 703 142
rect 637 17 703 108
rect 737 120 787 176
rect 737 86 753 120
rect 737 70 787 86
rect 823 210 889 226
rect 823 176 839 210
rect 873 176 889 210
rect 823 120 889 176
rect 823 86 839 120
rect 873 86 889 120
rect 823 17 889 86
rect 923 210 973 384
rect 1007 316 1018 350
rect 1052 316 1061 350
rect 1007 310 1061 316
rect 1007 276 1018 310
rect 1052 276 1061 310
rect 1007 260 1061 276
rect 923 176 939 210
rect 923 120 973 176
rect 923 86 939 120
rect 923 70 973 86
rect 1009 205 1059 221
rect 1009 171 1025 205
rect 1009 120 1059 171
rect 1009 86 1025 120
rect 1009 17 1059 86
rect 1102 210 1145 384
rect 1180 316 1196 350
rect 1230 316 1246 350
rect 1180 310 1246 316
rect 1180 276 1196 310
rect 1230 276 1246 310
rect 1180 260 1246 276
rect 1102 176 1111 210
rect 1102 120 1145 176
rect 1102 86 1111 120
rect 1102 70 1145 86
rect 1181 205 1247 221
rect 1181 171 1197 205
rect 1231 171 1247 205
rect 1181 120 1247 171
rect 1181 86 1197 120
rect 1231 86 1247 120
rect 1181 17 1247 86
rect 1284 210 1331 384
rect 1368 316 1384 350
rect 1418 316 1434 350
rect 1368 310 1434 316
rect 1368 276 1384 310
rect 1418 276 1434 310
rect 1368 260 1434 276
rect 1284 176 1297 210
rect 1284 120 1331 176
rect 1284 86 1297 120
rect 1284 70 1331 86
rect 1367 205 1433 221
rect 1367 171 1383 205
rect 1417 171 1433 205
rect 1367 120 1433 171
rect 1367 86 1383 120
rect 1417 86 1433 120
rect 1367 17 1433 86
rect 1468 210 1517 384
rect 1653 380 1664 404
rect 1698 384 1714 424
rect 1754 580 1799 649
rect 1788 546 1799 580
rect 1754 506 1799 546
rect 1788 472 1799 506
rect 1754 434 1799 472
rect 1788 400 1799 434
rect 1838 580 1904 596
rect 1838 546 1854 580
rect 1888 546 1904 580
rect 1838 497 1904 546
rect 1838 463 1854 497
rect 1888 463 1904 497
rect 1838 424 1904 463
rect 1838 404 1854 424
rect 1754 384 1799 400
rect 1698 380 1703 384
rect 1552 316 1567 350
rect 1601 316 1618 350
rect 1552 310 1618 316
rect 1552 276 1568 310
rect 1602 276 1618 310
rect 1552 260 1618 276
rect 1468 176 1483 210
rect 1468 120 1517 176
rect 1468 86 1483 120
rect 1468 70 1517 86
rect 1553 205 1619 221
rect 1553 171 1569 205
rect 1603 171 1619 205
rect 1553 120 1619 171
rect 1553 86 1569 120
rect 1603 86 1619 120
rect 1553 17 1619 86
rect 1653 210 1703 380
rect 1839 380 1854 404
rect 1888 384 1904 424
rect 1944 580 1991 649
rect 1978 546 1991 580
rect 1944 506 1991 546
rect 1978 472 1991 506
rect 1944 434 1991 472
rect 1978 400 1991 434
rect 2028 580 2094 596
rect 2028 546 2044 580
rect 2078 546 2094 580
rect 2028 497 2094 546
rect 2028 463 2044 497
rect 2078 463 2094 497
rect 2028 424 2094 463
rect 2028 404 2044 424
rect 1944 384 1991 400
rect 2025 384 2044 404
rect 2078 384 2094 424
rect 2134 580 2177 649
rect 2168 546 2177 580
rect 2134 506 2177 546
rect 2168 472 2177 506
rect 2134 434 2177 472
rect 2168 400 2177 434
rect 2218 580 2284 596
rect 2218 546 2234 580
rect 2268 546 2284 580
rect 2218 497 2284 546
rect 2218 463 2234 497
rect 2268 463 2284 497
rect 2218 424 2284 463
rect 2218 404 2234 424
rect 2134 384 2177 400
rect 1888 380 1889 384
rect 1737 316 1753 350
rect 1787 316 1803 350
rect 1737 310 1803 316
rect 1737 276 1753 310
rect 1787 276 1803 310
rect 1737 260 1803 276
rect 1653 176 1669 210
rect 1653 120 1703 176
rect 1653 86 1669 120
rect 1653 70 1703 86
rect 1739 205 1805 221
rect 1739 171 1755 205
rect 1789 171 1805 205
rect 1739 120 1805 171
rect 1739 86 1755 120
rect 1789 86 1805 120
rect 1739 17 1805 86
rect 1839 210 1889 380
rect 1923 316 1938 350
rect 1972 316 1989 350
rect 1923 310 1989 316
rect 1923 276 1939 310
rect 1973 276 1989 310
rect 1923 260 1989 276
rect 1839 176 1855 210
rect 1839 120 1889 176
rect 1839 86 1855 120
rect 1839 70 1889 86
rect 1925 205 1991 221
rect 1925 171 1941 205
rect 1975 171 1991 205
rect 1925 120 1991 171
rect 1925 86 1941 120
rect 1975 86 1991 120
rect 1925 17 1991 86
rect 2025 210 2075 384
rect 2211 380 2234 404
rect 2268 380 2284 424
rect 2211 358 2284 380
rect 2324 580 2374 649
rect 2358 546 2374 580
rect 2324 497 2374 546
rect 2358 463 2374 497
rect 2324 414 2374 463
rect 2358 380 2374 414
rect 2324 364 2374 380
rect 2109 316 2125 350
rect 2159 316 2175 350
rect 2109 310 2175 316
rect 2109 276 2125 310
rect 2159 276 2175 310
rect 2109 260 2175 276
rect 2025 176 2041 210
rect 2025 120 2075 176
rect 2025 86 2041 120
rect 2025 70 2075 86
rect 2111 205 2177 221
rect 2111 171 2127 205
rect 2161 171 2177 205
rect 2111 120 2177 171
rect 2111 86 2127 120
rect 2161 86 2177 120
rect 2111 17 2177 86
rect 2211 210 2277 358
rect 2211 176 2227 210
rect 2261 176 2277 210
rect 2211 120 2277 176
rect 2211 86 2227 120
rect 2261 86 2277 120
rect 2211 70 2277 86
rect 2311 210 2377 226
rect 2311 176 2327 210
rect 2361 176 2377 210
rect 2311 120 2377 176
rect 2311 86 2327 120
rect 2361 86 2377 120
rect 2311 17 2377 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 946 418 980 424
rect 946 390 978 418
rect 978 390 980 418
rect 1124 418 1158 424
rect 1124 390 1158 418
rect 1304 418 1338 424
rect 1304 390 1338 418
rect 1484 418 1518 424
rect 1484 390 1518 418
rect 1664 414 1698 424
rect 845 316 879 350
rect 1018 316 1052 350
rect 1196 316 1230 350
rect 1384 316 1418 350
rect 1664 390 1698 414
rect 1854 414 1888 424
rect 1567 316 1601 350
rect 1854 390 1888 414
rect 2044 418 2078 424
rect 2044 390 2078 418
rect 2234 414 2268 424
rect 1753 316 1787 350
rect 1938 316 1972 350
rect 2234 390 2268 414
rect 2125 316 2159 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 932 424 2280 430
rect 932 390 946 424
rect 980 390 1124 424
rect 1158 390 1304 424
rect 1338 390 1484 424
rect 1518 390 1664 424
rect 1698 390 1854 424
rect 1888 390 2044 424
rect 2078 390 2234 424
rect 2268 390 2280 424
rect 932 384 2280 390
rect 831 350 2171 356
rect 831 316 845 350
rect 879 316 1018 350
rect 1052 316 1196 350
rect 1230 316 1384 350
rect 1418 316 1567 350
rect 1601 316 1753 350
rect 1787 316 1938 350
rect 1972 316 2125 350
rect 2159 316 2171 350
rect 831 310 2171 316
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
rlabel comment s 0 0 0 0 4 bufinv_16
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nbase s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 932 384 2280 430 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 2400 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3312056
string GDS_START 3291936
<< end >>
