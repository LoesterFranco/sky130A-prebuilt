magic
tech sky130A
magscale 1 2
timestamp 1599588201
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 53 109 137
rect 175 53 205 137
rect 259 53 289 137
rect 343 53 373 137
rect 441 47 471 177
<< pmoshvt >>
rect 79 297 109 381
rect 175 297 205 381
rect 247 297 277 381
rect 343 297 373 381
rect 441 297 471 497
<< ndiff >>
rect 388 137 441 177
rect 27 117 79 137
rect 27 83 35 117
rect 69 83 79 117
rect 27 53 79 83
rect 109 111 175 137
rect 109 77 125 111
rect 159 77 175 111
rect 109 53 175 77
rect 205 97 259 137
rect 205 63 215 97
rect 249 63 259 97
rect 205 53 259 63
rect 289 111 343 137
rect 289 77 299 111
rect 333 77 343 111
rect 289 53 343 77
rect 373 97 441 137
rect 373 63 393 97
rect 427 63 441 97
rect 373 53 441 63
rect 388 47 441 53
rect 471 135 525 177
rect 471 101 481 135
rect 515 101 525 135
rect 471 47 525 101
<< pdiff >>
rect 388 485 441 497
rect 388 451 396 485
rect 430 451 441 485
rect 388 417 441 451
rect 388 383 396 417
rect 430 383 441 417
rect 388 381 441 383
rect 27 354 79 381
rect 27 320 35 354
rect 69 320 79 354
rect 27 297 79 320
rect 109 297 175 381
rect 205 297 247 381
rect 277 297 343 381
rect 373 297 441 381
rect 471 454 525 497
rect 471 420 481 454
rect 515 420 525 454
rect 471 386 525 420
rect 471 352 481 386
rect 515 352 525 386
rect 471 297 525 352
<< ndiffc >>
rect 35 83 69 117
rect 125 77 159 111
rect 215 63 249 97
rect 299 77 333 111
rect 393 63 427 97
rect 481 101 515 135
<< pdiffc >>
rect 396 451 430 485
rect 396 383 430 417
rect 35 320 69 354
rect 481 420 515 454
rect 481 352 515 386
<< poly >>
rect 441 497 471 523
rect 241 473 307 483
rect 241 439 257 473
rect 291 439 307 473
rect 241 429 307 439
rect 79 381 109 407
rect 175 381 205 407
rect 247 381 277 429
rect 343 381 373 407
rect 79 265 109 297
rect 175 265 205 297
rect 25 249 109 265
rect 25 215 35 249
rect 69 215 109 249
rect 25 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 79 137 109 199
rect 175 137 205 199
rect 247 182 277 297
rect 343 265 373 297
rect 441 265 471 297
rect 327 249 381 265
rect 327 215 337 249
rect 371 215 381 249
rect 327 199 381 215
rect 423 249 478 265
rect 423 215 433 249
rect 467 215 478 249
rect 423 199 478 215
rect 247 181 288 182
rect 247 152 289 181
rect 259 137 289 152
rect 343 137 373 199
rect 441 177 471 199
rect 79 27 109 53
rect 175 27 205 53
rect 259 27 289 53
rect 343 27 373 53
rect 441 21 471 47
<< polycont >>
rect 257 439 291 473
rect 35 215 69 249
rect 161 215 195 249
rect 337 215 371 249
rect 433 215 467 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 383 485 439 527
rect 18 473 349 483
rect 18 439 257 473
rect 291 439 349 473
rect 18 425 349 439
rect 383 451 396 485
rect 430 451 439 485
rect 383 417 439 451
rect 18 357 336 391
rect 383 383 396 417
rect 430 383 439 417
rect 383 367 439 383
rect 481 454 535 493
rect 515 420 535 454
rect 481 386 535 420
rect 18 354 82 357
rect 18 320 35 354
rect 69 320 82 354
rect 302 333 336 357
rect 515 352 535 386
rect 18 299 82 320
rect 18 249 88 265
rect 18 215 35 249
rect 69 215 88 249
rect 18 151 88 215
rect 122 249 264 323
rect 302 299 447 333
rect 481 299 535 352
rect 413 265 447 299
rect 122 215 161 249
rect 195 215 264 249
rect 122 199 264 215
rect 298 249 379 265
rect 298 215 337 249
rect 371 215 379 249
rect 298 199 379 215
rect 413 249 467 265
rect 413 215 433 249
rect 413 199 467 215
rect 413 165 447 199
rect 125 131 447 165
rect 501 152 535 299
rect 481 135 535 152
rect 19 83 35 117
rect 69 83 85 117
rect 19 17 85 83
rect 125 111 159 131
rect 299 111 333 131
rect 125 61 159 77
rect 199 63 215 97
rect 249 63 265 97
rect 199 17 265 63
rect 515 101 535 135
rect 299 61 333 77
rect 367 63 393 97
rect 427 63 443 97
rect 481 83 535 101
rect 367 17 443 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel corelocali s 214 221 248 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 306 221 340 255 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel corelocali s 490 357 524 391 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel corelocali s 122 221 156 255 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 214 425 248 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 122 425 156 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 122 289 156 323 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 30 425 64 459 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel corelocali s 214 289 248 323 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel corelocali s 30 153 64 187 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 or4_1
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1069060
string GDS_START 1063038
string path 0.000 0.000 2.760 0.000 
<< end >>
