magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1472 561
rect 111 425 161 527
rect 279 425 329 527
rect 635 427 685 527
rect 17 289 337 323
rect 971 359 1021 527
rect 1055 391 1105 493
rect 1139 433 1189 527
rect 1223 391 1273 493
rect 1055 357 1273 391
rect 1307 365 1357 527
rect 17 215 115 289
rect 161 215 269 255
rect 303 249 337 289
rect 1223 331 1273 357
rect 303 215 379 249
rect 695 289 993 323
rect 695 265 729 289
rect 663 215 729 265
rect 763 215 887 255
rect 921 215 993 289
rect 1223 283 1384 331
rect 1322 181 1384 283
rect 35 17 69 179
rect 371 17 405 111
rect 539 17 677 111
rect 811 17 845 111
rect 979 17 1013 179
rect 1047 145 1384 181
rect 1047 55 1113 145
rect 1147 17 1181 111
rect 1215 55 1281 145
rect 1315 17 1349 111
rect 0 -17 1472 17
<< obsli1 >>
rect 27 391 77 493
rect 195 391 245 493
rect 363 459 581 493
rect 363 391 413 459
rect 531 427 581 459
rect 719 459 937 493
rect 719 427 769 459
rect 27 357 413 391
rect 371 291 413 357
rect 447 393 497 425
rect 803 393 853 425
rect 447 323 524 393
rect 627 357 853 393
rect 887 357 937 459
rect 627 333 661 357
rect 447 289 490 323
rect 447 283 524 289
rect 591 299 661 333
rect 447 181 489 283
rect 591 249 629 299
rect 523 215 629 249
rect 1027 289 1046 323
rect 1080 289 1092 323
rect 1027 249 1092 289
rect 1027 215 1288 249
rect 591 181 629 215
rect 103 95 153 181
rect 187 147 505 181
rect 187 129 254 147
rect 103 51 337 95
rect 439 51 505 147
rect 591 145 945 181
rect 711 51 777 145
rect 879 51 945 145
<< obsli1c >>
rect 490 289 524 323
rect 1046 289 1080 323
<< metal1 >>
rect 0 496 1472 592
rect 0 -48 1472 48
<< obsm1 >>
rect 478 323 536 329
rect 478 289 490 323
rect 524 320 536 323
rect 1034 323 1092 329
rect 1034 320 1046 323
rect 524 292 1046 320
rect 524 289 536 292
rect 478 283 536 289
rect 1034 289 1046 292
rect 1080 289 1092 323
rect 1034 283 1092 289
<< labels >>
rlabel locali s 921 215 993 289 6 A1_N
port 1 nsew signal input
rlabel locali s 695 289 993 323 6 A1_N
port 1 nsew signal input
rlabel locali s 695 265 729 289 6 A1_N
port 1 nsew signal input
rlabel locali s 663 215 729 265 6 A1_N
port 1 nsew signal input
rlabel locali s 763 215 887 255 6 A2_N
port 2 nsew signal input
rlabel locali s 303 249 337 289 6 B1
port 3 nsew signal input
rlabel locali s 303 215 379 249 6 B1
port 3 nsew signal input
rlabel locali s 17 289 337 323 6 B1
port 3 nsew signal input
rlabel locali s 17 215 115 289 6 B1
port 3 nsew signal input
rlabel locali s 161 215 269 255 6 B2
port 4 nsew signal input
rlabel locali s 1322 181 1384 283 6 X
port 5 nsew signal output
rlabel locali s 1223 391 1273 493 6 X
port 5 nsew signal output
rlabel locali s 1223 331 1273 357 6 X
port 5 nsew signal output
rlabel locali s 1223 283 1384 331 6 X
port 5 nsew signal output
rlabel locali s 1215 55 1281 145 6 X
port 5 nsew signal output
rlabel locali s 1055 391 1105 493 6 X
port 5 nsew signal output
rlabel locali s 1055 357 1273 391 6 X
port 5 nsew signal output
rlabel locali s 1047 145 1384 181 6 X
port 5 nsew signal output
rlabel locali s 1047 55 1113 145 6 X
port 5 nsew signal output
rlabel locali s 1315 17 1349 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1147 17 1181 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 979 17 1013 179 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 811 17 845 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 539 17 677 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 371 17 405 111 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 35 17 69 179 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 1307 365 1357 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1139 433 1189 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 971 359 1021 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 635 427 685 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 279 425 329 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 111 425 161 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3475012
string GDS_START 3463608
<< end >>
