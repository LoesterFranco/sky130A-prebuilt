magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 84 47 114 177
rect 180 47 210 177
rect 276 47 306 177
rect 372 47 402 177
rect 575 47 605 177
rect 679 47 709 177
rect 771 47 801 177
rect 857 47 887 177
rect 961 47 991 177
rect 1045 47 1075 177
<< pmoshvt >>
rect 86 297 122 497
rect 182 297 218 497
rect 278 297 314 497
rect 374 297 410 497
rect 577 297 613 497
rect 671 297 707 497
rect 765 297 801 497
rect 859 297 895 497
rect 953 297 989 497
rect 1047 297 1083 497
<< ndiff >>
rect 27 89 84 177
rect 27 55 39 89
rect 73 55 84 89
rect 27 47 84 55
rect 114 157 180 177
rect 114 123 135 157
rect 169 123 180 157
rect 114 47 180 123
rect 210 89 276 177
rect 210 55 231 89
rect 265 55 276 89
rect 210 47 276 55
rect 306 157 372 177
rect 306 123 327 157
rect 361 123 372 157
rect 306 47 372 123
rect 402 89 575 177
rect 402 55 445 89
rect 479 55 527 89
rect 561 55 575 89
rect 402 47 575 55
rect 605 169 679 177
rect 605 135 625 169
rect 659 135 679 169
rect 605 101 679 135
rect 605 67 625 101
rect 659 67 679 101
rect 605 47 679 67
rect 709 89 771 177
rect 709 55 727 89
rect 761 55 771 89
rect 709 47 771 55
rect 801 47 857 177
rect 887 131 961 177
rect 887 97 907 131
rect 941 97 961 131
rect 887 47 961 97
rect 991 47 1045 177
rect 1075 161 1137 177
rect 1075 127 1095 161
rect 1129 127 1137 161
rect 1075 93 1137 127
rect 1075 59 1095 93
rect 1129 59 1137 93
rect 1075 47 1137 59
<< pdiff >>
rect 27 489 86 497
rect 27 455 39 489
rect 73 455 86 489
rect 27 421 86 455
rect 27 387 39 421
rect 73 387 86 421
rect 27 297 86 387
rect 122 421 182 497
rect 122 387 135 421
rect 169 387 182 421
rect 122 351 182 387
rect 122 317 135 351
rect 169 317 182 351
rect 122 297 182 317
rect 218 489 278 497
rect 218 455 231 489
rect 265 455 278 489
rect 218 421 278 455
rect 218 387 231 421
rect 265 387 278 421
rect 218 297 278 387
rect 314 421 374 497
rect 314 387 327 421
rect 361 387 374 421
rect 314 351 374 387
rect 314 317 327 351
rect 361 317 374 351
rect 314 297 374 317
rect 410 489 469 497
rect 410 455 423 489
rect 457 455 469 489
rect 410 421 469 455
rect 410 387 423 421
rect 457 387 469 421
rect 410 353 469 387
rect 410 319 423 353
rect 457 319 469 353
rect 410 297 469 319
rect 523 459 577 497
rect 523 425 531 459
rect 565 425 577 459
rect 523 389 577 425
rect 523 355 531 389
rect 565 355 577 389
rect 523 297 577 355
rect 613 409 671 497
rect 613 375 625 409
rect 659 375 671 409
rect 613 341 671 375
rect 613 307 625 341
rect 659 307 671 341
rect 613 297 671 307
rect 707 428 765 497
rect 707 394 719 428
rect 753 394 765 428
rect 707 339 765 394
rect 707 305 719 339
rect 753 305 765 339
rect 707 297 765 305
rect 801 489 859 497
rect 801 455 813 489
rect 847 455 859 489
rect 801 297 859 455
rect 895 477 953 497
rect 895 443 907 477
rect 941 443 953 477
rect 895 404 953 443
rect 895 370 907 404
rect 941 370 953 404
rect 895 297 953 370
rect 989 489 1047 497
rect 989 455 1001 489
rect 1035 455 1047 489
rect 989 297 1047 455
rect 1083 479 1164 497
rect 1083 445 1122 479
rect 1156 445 1164 479
rect 1083 411 1164 445
rect 1083 377 1122 411
rect 1156 377 1164 411
rect 1083 343 1164 377
rect 1083 309 1122 343
rect 1156 309 1164 343
rect 1083 297 1164 309
<< ndiffc >>
rect 39 55 73 89
rect 135 123 169 157
rect 231 55 265 89
rect 327 123 361 157
rect 445 55 479 89
rect 527 55 561 89
rect 625 135 659 169
rect 625 67 659 101
rect 727 55 761 89
rect 907 97 941 131
rect 1095 127 1129 161
rect 1095 59 1129 93
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 135 387 169 421
rect 135 317 169 351
rect 231 455 265 489
rect 231 387 265 421
rect 327 387 361 421
rect 327 317 361 351
rect 423 455 457 489
rect 423 387 457 421
rect 423 319 457 353
rect 531 425 565 459
rect 531 355 565 389
rect 625 375 659 409
rect 625 307 659 341
rect 719 394 753 428
rect 719 305 753 339
rect 813 455 847 489
rect 907 443 941 477
rect 907 370 941 404
rect 1001 455 1035 489
rect 1122 445 1156 479
rect 1122 377 1156 411
rect 1122 309 1156 343
<< poly >>
rect 86 497 122 523
rect 182 497 218 523
rect 278 497 314 523
rect 374 497 410 523
rect 577 497 613 523
rect 671 497 707 523
rect 765 497 801 523
rect 859 497 895 523
rect 953 497 989 523
rect 1047 497 1083 523
rect 86 282 122 297
rect 182 282 218 297
rect 278 282 314 297
rect 374 282 410 297
rect 577 282 613 297
rect 671 282 707 297
rect 765 282 801 297
rect 859 282 895 297
rect 953 282 989 297
rect 1047 282 1083 297
rect 84 265 124 282
rect 180 265 220 282
rect 276 265 316 282
rect 372 265 412 282
rect 575 265 615 282
rect 669 265 709 282
rect 763 265 803 282
rect 857 265 897 282
rect 951 265 991 282
rect 84 249 435 265
rect 84 215 235 249
rect 269 215 303 249
rect 337 215 381 249
rect 415 215 435 249
rect 84 199 435 215
rect 537 249 709 265
rect 537 215 547 249
rect 581 215 709 249
rect 537 199 709 215
rect 751 249 815 265
rect 751 215 761 249
rect 795 215 815 249
rect 751 199 815 215
rect 857 249 991 265
rect 857 215 901 249
rect 935 215 991 249
rect 857 199 991 215
rect 84 177 114 199
rect 180 177 210 199
rect 276 177 306 199
rect 372 177 402 199
rect 575 177 605 199
rect 679 177 709 199
rect 771 177 801 199
rect 857 177 887 199
rect 961 177 991 199
rect 1045 265 1085 282
rect 1045 249 1109 265
rect 1045 215 1055 249
rect 1089 215 1109 249
rect 1045 199 1109 215
rect 1045 177 1075 199
rect 84 21 114 47
rect 180 21 210 47
rect 276 21 306 47
rect 372 21 402 47
rect 575 21 605 47
rect 679 21 709 47
rect 771 21 801 47
rect 857 21 887 47
rect 961 21 991 47
rect 1045 21 1075 47
<< polycont >>
rect 235 215 269 249
rect 303 215 337 249
rect 381 215 415 249
rect 547 215 581 249
rect 761 215 795 249
rect 901 215 935 249
rect 1055 215 1089 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 23 489 89 527
rect 23 455 39 489
rect 73 455 89 489
rect 23 421 89 455
rect 205 489 281 527
rect 205 455 231 489
rect 265 455 281 489
rect 23 387 39 421
rect 73 387 89 421
rect 135 421 169 437
rect 205 421 281 455
rect 413 489 463 527
rect 413 455 423 489
rect 457 455 463 489
rect 205 387 231 421
rect 265 387 281 421
rect 327 421 377 437
rect 361 387 377 421
rect 135 351 169 387
rect 327 351 377 387
rect 29 317 135 351
rect 169 317 327 351
rect 361 317 377 351
rect 413 421 463 455
rect 413 387 423 421
rect 457 387 463 421
rect 413 353 463 387
rect 413 319 423 353
rect 457 319 463 353
rect 531 459 753 493
rect 717 428 753 459
rect 787 489 863 527
rect 787 455 813 489
rect 847 455 863 489
rect 907 477 941 493
rect 531 389 565 425
rect 531 339 565 355
rect 625 409 659 425
rect 625 341 659 375
rect 29 157 136 317
rect 413 303 463 319
rect 170 249 460 265
rect 170 215 235 249
rect 269 215 303 249
rect 337 215 381 249
rect 415 215 460 249
rect 170 199 460 215
rect 500 249 581 305
rect 500 215 547 249
rect 500 199 581 215
rect 426 157 460 199
rect 625 169 659 307
rect 717 394 719 428
rect 975 489 1051 527
rect 975 455 1001 489
rect 1035 455 1051 489
rect 907 404 941 443
rect 1106 445 1122 479
rect 1156 445 1172 479
rect 1106 411 1172 445
rect 1106 404 1122 411
rect 753 394 907 404
rect 717 370 907 394
rect 941 377 1122 404
rect 1156 377 1172 411
rect 941 370 1172 377
rect 717 339 753 370
rect 717 305 719 339
rect 1121 343 1172 370
rect 717 289 753 305
rect 789 302 1087 336
rect 789 255 834 302
rect 1027 258 1087 302
rect 1121 309 1122 343
rect 1156 309 1172 343
rect 1121 292 1172 309
rect 745 249 834 255
rect 745 215 761 249
rect 795 215 834 249
rect 745 202 834 215
rect 868 249 993 255
rect 868 215 901 249
rect 935 215 993 249
rect 868 202 993 215
rect 1027 249 1120 258
rect 1027 215 1055 249
rect 1089 215 1120 249
rect 1027 211 1120 215
rect 29 123 135 157
rect 169 123 327 157
rect 361 123 377 157
rect 426 135 625 157
rect 659 135 953 168
rect 426 134 953 135
rect 426 123 659 134
rect 625 101 659 123
rect 21 55 39 89
rect 73 55 89 89
rect 21 17 89 55
rect 205 55 231 89
rect 265 55 281 89
rect 205 17 281 55
rect 422 55 445 89
rect 479 55 527 89
rect 561 55 577 89
rect 422 17 577 55
rect 897 131 953 134
rect 897 97 907 131
rect 941 97 953 131
rect 625 51 659 67
rect 711 55 727 89
rect 761 55 777 89
rect 897 81 953 97
rect 1089 161 1145 177
rect 1089 127 1095 161
rect 1129 127 1145 161
rect 1089 93 1145 127
rect 711 17 777 55
rect 1089 59 1095 93
rect 1129 59 1145 93
rect 1089 17 1145 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel corelocali s 970 306 970 306 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 878 238 878 238 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 29 289 63 323 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 510 238 510 238 0 FreeSans 340 0 0 0 B1
port 3 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1194602
string GDS_START 1186030
<< end >>
