magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< locali >>
rect 21 260 87 356
rect 121 252 228 356
rect 339 364 488 440
rect 339 184 405 364
rect 585 270 651 430
rect 693 270 759 356
rect 793 270 889 356
rect 937 270 1031 356
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 440 73 596
rect 113 508 179 596
rect 315 542 381 649
rect 529 542 595 649
rect 653 581 933 615
rect 653 542 726 581
rect 767 508 833 547
rect 113 474 833 508
rect 23 390 305 440
rect 271 218 305 390
rect 23 184 305 218
rect 446 236 512 318
rect 767 390 833 474
rect 867 390 933 581
rect 967 390 1033 649
rect 446 202 750 236
rect 23 78 73 184
rect 271 150 305 184
rect 446 150 480 202
rect 187 17 237 150
rect 271 116 480 150
rect 553 104 619 168
rect 653 140 750 202
rect 784 202 1028 236
rect 784 104 818 202
rect 441 17 507 82
rect 553 70 818 104
rect 852 17 918 168
rect 962 70 1028 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel locali s 585 270 651 430 6 A1
port 1 nsew signal input
rlabel locali s 937 270 1031 356 6 A2
port 2 nsew signal input
rlabel locali s 693 270 759 356 6 B1
port 3 nsew signal input
rlabel locali s 793 270 889 356 6 B2
port 4 nsew signal input
rlabel locali s 21 260 87 356 6 C1
port 5 nsew signal input
rlabel locali s 121 252 228 356 6 C2
port 6 nsew signal input
rlabel locali s 339 364 488 440 6 X
port 7 nsew signal output
rlabel locali s 339 184 405 364 6 X
port 7 nsew signal output
rlabel metal1 s 0 -49 1056 49 8 VGND
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1056 715 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3493034
string GDS_START 3484380
<< end >>
