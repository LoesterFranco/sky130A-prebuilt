magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 24 153 85 361
rect 305 157 373 423
rect 460 299 817 335
rect 460 249 535 299
rect 459 215 535 249
rect 571 199 713 265
rect 747 199 817 299
rect 305 123 672 157
rect 305 51 374 123
rect 596 51 672 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 19 416 85 527
rect 220 457 483 493
rect 129 257 165 453
rect 220 359 270 457
rect 129 214 271 257
rect 129 106 165 214
rect 53 72 165 106
rect 217 17 265 177
rect 407 405 483 457
rect 527 439 561 527
rect 622 421 656 493
rect 692 455 768 527
rect 812 421 864 493
rect 622 405 864 421
rect 407 371 864 405
rect 428 17 494 89
rect 798 17 866 157
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 571 199 713 265 6 A1
port 1 nsew signal input
rlabel locali s 747 199 817 299 6 A2
port 2 nsew signal input
rlabel locali s 460 299 817 335 6 A2
port 2 nsew signal input
rlabel locali s 460 249 535 299 6 A2
port 2 nsew signal input
rlabel locali s 459 215 535 249 6 A2
port 2 nsew signal input
rlabel locali s 24 153 85 361 6 B1_N
port 3 nsew signal input
rlabel locali s 596 51 672 123 6 Y
port 4 nsew signal output
rlabel locali s 305 157 373 423 6 Y
port 4 nsew signal output
rlabel locali s 305 123 672 157 6 Y
port 4 nsew signal output
rlabel locali s 305 51 374 123 6 Y
port 4 nsew signal output
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1163918
string GDS_START 1156918
<< end >>
