magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 2024 561
rect 35 289 69 527
rect 203 367 237 527
rect 371 367 405 527
rect 539 367 573 527
rect 607 323 673 493
rect 707 367 741 527
rect 775 323 841 493
rect 875 367 909 527
rect 943 323 1009 493
rect 1043 367 1077 527
rect 1111 323 1177 493
rect 1211 367 1245 527
rect 1279 323 1345 493
rect 1379 367 1413 527
rect 1447 323 1513 493
rect 1547 367 1581 527
rect 1615 323 1681 493
rect 1715 367 1749 527
rect 1783 323 1849 493
rect 1883 367 1917 527
rect 1952 323 2007 472
rect 607 289 2007 323
rect 17 215 497 255
rect 1931 181 2007 289
rect 35 17 69 181
rect 607 147 2007 181
rect 203 17 237 113
rect 371 17 405 113
rect 539 17 573 113
rect 607 52 673 147
rect 607 51 657 52
rect 707 17 741 113
rect 775 52 841 147
rect 791 51 825 52
rect 875 17 909 113
rect 943 52 1009 147
rect 959 51 993 52
rect 1043 17 1077 113
rect 1111 52 1177 147
rect 1211 17 1245 113
rect 1279 52 1345 147
rect 1379 17 1413 113
rect 1447 52 1513 147
rect 1547 17 1581 113
rect 1615 52 1681 147
rect 1715 17 1749 113
rect 1783 52 1849 147
rect 1883 17 1917 113
rect 1952 73 2007 147
rect 0 -17 2024 17
<< obsli1 >>
rect 103 323 169 493
rect 271 323 337 493
rect 439 323 505 493
rect 103 289 573 323
rect 538 255 573 289
rect 538 215 1882 255
rect 538 181 573 215
rect 103 147 573 181
rect 103 52 169 147
rect 271 52 337 147
rect 439 52 505 147
<< metal1 >>
rect 0 496 2024 592
rect 0 -48 2024 48
<< labels >>
rlabel locali s 17 215 497 255 6 A
port 1 nsew signal input
rlabel locali s 1952 323 2007 472 6 X
port 2 nsew signal output
rlabel locali s 1952 73 2007 147 6 X
port 2 nsew signal output
rlabel locali s 1931 181 2007 289 6 X
port 2 nsew signal output
rlabel locali s 1783 323 1849 493 6 X
port 2 nsew signal output
rlabel locali s 1783 52 1849 147 6 X
port 2 nsew signal output
rlabel locali s 1615 323 1681 493 6 X
port 2 nsew signal output
rlabel locali s 1615 52 1681 147 6 X
port 2 nsew signal output
rlabel locali s 1447 323 1513 493 6 X
port 2 nsew signal output
rlabel locali s 1447 52 1513 147 6 X
port 2 nsew signal output
rlabel locali s 1279 323 1345 493 6 X
port 2 nsew signal output
rlabel locali s 1279 52 1345 147 6 X
port 2 nsew signal output
rlabel locali s 1111 323 1177 493 6 X
port 2 nsew signal output
rlabel locali s 1111 52 1177 147 6 X
port 2 nsew signal output
rlabel locali s 959 51 993 52 6 X
port 2 nsew signal output
rlabel locali s 943 323 1009 493 6 X
port 2 nsew signal output
rlabel locali s 943 52 1009 147 6 X
port 2 nsew signal output
rlabel locali s 791 51 825 52 6 X
port 2 nsew signal output
rlabel locali s 775 323 841 493 6 X
port 2 nsew signal output
rlabel locali s 775 52 841 147 6 X
port 2 nsew signal output
rlabel locali s 607 323 673 493 6 X
port 2 nsew signal output
rlabel locali s 607 289 2007 323 6 X
port 2 nsew signal output
rlabel locali s 607 147 2007 181 6 X
port 2 nsew signal output
rlabel locali s 607 52 673 147 6 X
port 2 nsew signal output
rlabel locali s 607 51 657 52 6 X
port 2 nsew signal output
rlabel locali s 1883 17 1917 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1715 17 1749 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1547 17 1581 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1379 17 1413 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1211 17 1245 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1043 17 1077 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 875 17 909 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 707 17 741 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 539 17 573 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 371 17 405 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 203 17 237 113 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 35 17 69 181 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2024 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1883 367 1917 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1715 367 1749 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1547 367 1581 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1379 367 1413 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1211 367 1245 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1043 367 1077 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 875 367 909 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 707 367 741 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 539 367 573 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 371 367 405 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 203 367 237 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 35 289 69 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 2024 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3031450
string GDS_START 3015974
<< end >>
