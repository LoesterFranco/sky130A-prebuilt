magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 25 260 99 356
rect 391 236 551 302
rect 2143 270 2223 356
rect 2329 404 2363 596
rect 2329 370 2397 404
rect 2363 236 2397 370
rect 2703 388 2769 596
rect 2703 354 2807 388
rect 2326 88 2397 236
rect 2773 220 2807 354
rect 2708 170 2807 220
rect 2708 70 2760 170
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 21 424 87 596
rect 127 458 161 649
rect 201 581 425 615
rect 21 390 167 424
rect 133 326 167 390
rect 201 364 289 581
rect 133 260 221 326
rect 133 226 167 260
rect 255 226 289 364
rect 23 192 167 226
rect 23 70 73 192
rect 109 17 175 158
rect 211 70 289 226
rect 323 202 357 547
rect 391 371 425 581
rect 459 505 493 649
rect 527 581 921 615
rect 527 471 561 581
rect 617 513 714 547
rect 473 405 561 471
rect 595 371 646 471
rect 391 337 646 371
rect 601 291 646 337
rect 680 359 714 513
rect 748 427 798 547
rect 837 498 921 581
rect 1011 532 1077 649
rect 1113 498 1179 596
rect 1219 532 1285 649
rect 837 464 1276 498
rect 837 461 955 464
rect 748 393 887 427
rect 680 325 819 359
rect 743 293 819 325
rect 601 276 709 291
rect 601 242 607 276
rect 641 242 709 276
rect 601 225 709 242
rect 323 168 556 202
rect 743 191 777 293
rect 853 259 887 393
rect 323 115 373 168
rect 409 17 488 134
rect 522 85 556 168
rect 596 157 777 191
rect 811 225 887 259
rect 921 259 955 461
rect 1083 424 1149 430
rect 1083 390 1087 424
rect 1121 390 1149 424
rect 989 322 1049 388
rect 1083 326 1149 390
rect 1210 326 1276 464
rect 1393 420 1491 596
rect 1602 594 1668 649
rect 1714 560 1780 596
rect 1821 594 1887 649
rect 2012 560 2078 596
rect 1015 292 1049 322
rect 921 225 981 259
rect 1015 258 1283 292
rect 596 119 662 157
rect 811 123 845 225
rect 947 224 981 225
rect 698 85 845 123
rect 522 51 845 85
rect 879 87 913 191
rect 947 121 1015 224
rect 1049 87 1115 205
rect 879 53 1115 87
rect 1149 17 1215 205
rect 1249 102 1283 258
rect 1357 282 1423 382
rect 1457 378 1491 420
rect 1585 526 2078 560
rect 2223 526 2289 649
rect 1585 412 1651 526
rect 2012 492 2078 526
rect 1685 458 1978 492
rect 2012 458 2292 492
rect 1685 378 1719 458
rect 1457 344 1719 378
rect 1753 390 1759 424
rect 1793 390 1799 424
rect 1753 356 1799 390
rect 1944 378 1978 458
rect 2075 390 2184 424
rect 1537 282 1587 310
rect 1357 276 1587 282
rect 1357 242 1375 276
rect 1409 242 1587 276
rect 1357 236 1587 242
rect 1621 202 1655 344
rect 1753 290 1832 356
rect 1944 344 2041 378
rect 1874 236 1940 310
rect 1982 294 2041 344
rect 2075 236 2109 390
rect 2258 336 2292 458
rect 2403 438 2469 649
rect 2258 270 2329 336
rect 1330 136 1655 202
rect 1689 202 2198 236
rect 1689 102 1723 202
rect 2258 168 2292 270
rect 2509 364 2575 572
rect 2613 364 2663 649
rect 2809 422 2859 649
rect 2527 320 2575 364
rect 2527 254 2739 320
rect 1249 68 1723 102
rect 1757 17 1791 168
rect 1827 85 1877 168
rect 1921 134 2292 168
rect 1921 119 1987 134
rect 2022 85 2088 100
rect 1827 51 2088 85
rect 2133 17 2290 100
rect 2431 17 2481 252
rect 2527 70 2577 254
rect 2619 17 2674 210
rect 2794 17 2860 136
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 607 242 641 276
rect 1087 390 1121 424
rect 1759 390 1793 424
rect 1375 242 1409 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 0 616 50 617
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1121 393 1759 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 0 49 50 50
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< obsm1 >>
rect 595 276 653 282
rect 595 242 607 276
rect 641 273 653 276
rect 1363 276 1421 282
rect 1363 273 1375 276
rect 641 245 1375 273
rect 641 242 653 245
rect 595 236 653 242
rect 1363 242 1375 245
rect 1409 242 1421 276
rect 1363 236 1421 242
<< labels >>
rlabel locali s 391 236 551 302 6 D
port 1 nsew signal input
rlabel locali s 2773 220 2807 354 6 Q
port 2 nsew signal output
rlabel locali s 2708 170 2807 220 6 Q
port 2 nsew signal output
rlabel locali s 2708 70 2760 170 6 Q
port 2 nsew signal output
rlabel locali s 2703 388 2769 596 6 Q
port 2 nsew signal output
rlabel locali s 2703 354 2807 388 6 Q
port 2 nsew signal output
rlabel locali s 2363 236 2397 370 6 Q_N
port 3 nsew signal output
rlabel locali s 2329 404 2363 596 6 Q_N
port 3 nsew signal output
rlabel locali s 2329 370 2397 404 6 Q_N
port 3 nsew signal output
rlabel locali s 2326 88 2397 236 6 Q_N
port 3 nsew signal output
rlabel locali s 2143 270 2223 356 6 RESET_B
port 4 nsew signal input
rlabel metal1 s 1747 421 1805 430 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1747 384 1805 393 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1075 421 1133 430 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1075 393 1805 421 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1075 384 1133 393 6 SET_B
port 5 nsew signal input
rlabel locali s 25 260 99 356 6 CLK_N
port 6 nsew clock input
rlabel metal1 s 0 -49 2880 49 8 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 617 2880 715 6 VPWR
port 10 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2753466
string GDS_START 2732014
<< end >>
