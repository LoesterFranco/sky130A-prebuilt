magic
tech sky130A
magscale 1 2
timestamp 1599588214
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 0 0 1728 49
<< scnmos >>
rect 92 81 122 209
rect 194 81 224 209
rect 299 81 329 209
rect 397 169 427 253
rect 499 125 529 253
rect 599 125 629 253
rect 813 89 843 237
rect 1027 74 1057 202
rect 1127 74 1157 202
rect 1339 162 1369 246
rect 1528 98 1558 246
rect 1614 98 1644 246
<< pmoshvt >>
rect 86 373 116 573
rect 194 373 224 573
rect 302 373 332 541
rect 424 373 454 501
rect 518 373 548 501
rect 626 373 656 541
rect 848 368 878 592
rect 1064 399 1094 567
rect 1187 399 1217 567
rect 1387 368 1417 496
rect 1523 368 1553 592
rect 1613 368 1643 592
<< ndiff >>
rect 347 209 397 253
rect 35 197 92 209
rect 35 163 47 197
rect 81 163 92 197
rect 35 127 92 163
rect 35 93 47 127
rect 81 93 92 127
rect 35 81 92 93
rect 122 173 194 209
rect 122 139 133 173
rect 167 139 194 173
rect 122 81 194 139
rect 224 197 299 209
rect 224 163 235 197
rect 269 163 299 197
rect 224 127 299 163
rect 224 93 235 127
rect 269 93 299 127
rect 224 81 299 93
rect 329 177 397 209
rect 329 143 340 177
rect 374 169 397 177
rect 427 239 499 253
rect 427 205 438 239
rect 472 205 499 239
rect 427 169 499 205
rect 374 143 382 169
rect 329 81 382 143
rect 449 125 499 169
rect 529 241 599 253
rect 529 207 543 241
rect 577 207 599 241
rect 529 125 599 207
rect 629 125 702 253
rect 644 89 702 125
rect 756 225 813 237
rect 756 191 768 225
rect 802 191 813 225
rect 756 89 813 191
rect 843 89 916 237
rect 1282 234 1339 246
rect 644 55 656 89
rect 690 55 702 89
rect 644 43 702 55
rect 858 55 870 89
rect 904 55 916 89
rect 970 193 1027 202
rect 970 159 982 193
rect 1016 159 1027 193
rect 970 120 1027 159
rect 970 86 982 120
rect 1016 86 1027 120
rect 970 74 1027 86
rect 1057 193 1127 202
rect 1057 159 1082 193
rect 1116 159 1127 193
rect 1057 116 1127 159
rect 1057 82 1082 116
rect 1116 82 1127 116
rect 1057 74 1127 82
rect 1157 179 1228 202
rect 1157 145 1182 179
rect 1216 145 1228 179
rect 1282 200 1294 234
rect 1328 200 1339 234
rect 1282 162 1339 200
rect 1369 168 1528 246
rect 1369 162 1462 168
rect 1157 74 1228 145
rect 1384 134 1462 162
rect 1496 134 1528 168
rect 1384 98 1528 134
rect 1558 218 1614 246
rect 1558 184 1569 218
rect 1603 184 1614 218
rect 1558 144 1614 184
rect 1558 110 1569 144
rect 1603 110 1614 144
rect 1558 98 1614 110
rect 1644 234 1701 246
rect 1644 200 1655 234
rect 1689 200 1701 234
rect 1644 144 1701 200
rect 1644 110 1655 144
rect 1689 110 1701 144
rect 1644 98 1701 110
rect 1384 82 1513 98
rect 858 43 916 55
rect 1384 48 1396 82
rect 1430 48 1467 82
rect 1501 48 1513 82
rect 1384 36 1513 48
<< pdiff >>
rect 27 561 86 573
rect 27 527 39 561
rect 73 527 86 561
rect 27 492 86 527
rect 27 458 39 492
rect 73 458 86 492
rect 27 373 86 458
rect 116 521 194 573
rect 116 487 132 521
rect 166 487 194 521
rect 116 373 194 487
rect 224 561 281 573
rect 224 527 239 561
rect 273 541 281 561
rect 273 527 302 541
rect 224 440 302 527
rect 224 406 239 440
rect 273 406 302 440
rect 224 373 302 406
rect 332 501 386 541
rect 674 576 730 588
rect 674 542 685 576
rect 719 542 730 576
rect 674 541 730 542
rect 567 508 626 541
rect 567 501 579 508
rect 332 441 424 501
rect 332 407 377 441
rect 411 407 424 441
rect 332 373 424 407
rect 454 489 518 501
rect 454 455 471 489
rect 505 455 518 489
rect 454 419 518 455
rect 454 385 471 419
rect 505 385 518 419
rect 454 373 518 385
rect 548 474 579 501
rect 613 474 626 508
rect 548 425 626 474
rect 548 391 579 425
rect 613 391 626 425
rect 548 373 626 391
rect 656 373 730 541
rect 896 597 952 609
rect 896 592 907 597
rect 790 440 848 592
rect 790 406 801 440
rect 835 406 848 440
rect 790 368 848 406
rect 878 563 907 592
rect 941 563 952 597
rect 1112 581 1169 593
rect 1112 567 1123 581
rect 878 368 952 563
rect 1006 445 1064 567
rect 1006 411 1017 445
rect 1051 411 1064 445
rect 1006 399 1064 411
rect 1094 547 1123 567
rect 1157 567 1169 581
rect 1464 580 1523 592
rect 1157 547 1187 567
rect 1094 399 1187 547
rect 1217 531 1275 567
rect 1217 497 1230 531
rect 1264 497 1275 531
rect 1464 546 1476 580
rect 1510 546 1523 580
rect 1217 445 1275 497
rect 1464 508 1523 546
rect 1464 496 1476 508
rect 1217 411 1230 445
rect 1264 411 1275 445
rect 1217 399 1275 411
rect 1329 462 1387 496
rect 1329 428 1340 462
rect 1374 428 1387 462
rect 1329 368 1387 428
rect 1417 474 1476 496
rect 1510 474 1523 508
rect 1417 368 1523 474
rect 1553 580 1613 592
rect 1553 546 1566 580
rect 1600 546 1613 580
rect 1553 499 1613 546
rect 1553 465 1566 499
rect 1600 465 1613 499
rect 1553 418 1613 465
rect 1553 384 1566 418
rect 1600 384 1613 418
rect 1553 368 1613 384
rect 1643 580 1701 592
rect 1643 546 1656 580
rect 1690 546 1701 580
rect 1643 497 1701 546
rect 1643 463 1656 497
rect 1690 463 1701 497
rect 1643 414 1701 463
rect 1643 380 1656 414
rect 1690 380 1701 414
rect 1643 368 1701 380
<< ndiffc >>
rect 47 163 81 197
rect 47 93 81 127
rect 133 139 167 173
rect 235 163 269 197
rect 235 93 269 127
rect 340 143 374 177
rect 438 205 472 239
rect 543 207 577 241
rect 768 191 802 225
rect 656 55 690 89
rect 870 55 904 89
rect 982 159 1016 193
rect 982 86 1016 120
rect 1082 159 1116 193
rect 1082 82 1116 116
rect 1182 145 1216 179
rect 1294 200 1328 234
rect 1462 134 1496 168
rect 1569 184 1603 218
rect 1569 110 1603 144
rect 1655 200 1689 234
rect 1655 110 1689 144
rect 1396 48 1430 82
rect 1467 48 1501 82
<< pdiffc >>
rect 39 527 73 561
rect 39 458 73 492
rect 132 487 166 521
rect 239 527 273 561
rect 239 406 273 440
rect 685 542 719 576
rect 377 407 411 441
rect 471 455 505 489
rect 471 385 505 419
rect 579 474 613 508
rect 579 391 613 425
rect 801 406 835 440
rect 907 563 941 597
rect 1017 411 1051 445
rect 1123 547 1157 581
rect 1230 497 1264 531
rect 1476 546 1510 580
rect 1230 411 1264 445
rect 1340 428 1374 462
rect 1476 474 1510 508
rect 1566 546 1600 580
rect 1566 465 1600 499
rect 1566 384 1600 418
rect 1656 546 1690 580
rect 1656 463 1690 497
rect 1656 380 1690 414
<< poly >>
rect 299 615 775 645
rect 86 573 116 599
rect 194 573 224 599
rect 299 556 335 615
rect 302 541 332 556
rect 424 501 454 527
rect 515 516 551 615
rect 626 541 656 567
rect 518 501 548 516
rect 86 358 116 373
rect 194 358 224 373
rect 302 358 332 373
rect 424 358 454 373
rect 518 358 548 373
rect 626 358 656 373
rect 83 313 119 358
rect 191 341 227 358
rect 191 325 257 341
rect 83 297 149 313
rect 83 263 99 297
rect 133 263 149 297
rect 191 291 207 325
rect 241 291 257 325
rect 191 275 257 291
rect 299 301 335 358
rect 83 247 149 263
rect 92 209 122 247
rect 194 209 224 275
rect 299 209 329 301
rect 421 298 457 358
rect 515 331 551 358
rect 623 341 659 358
rect 397 268 457 298
rect 499 301 551 331
rect 599 325 697 341
rect 397 253 427 268
rect 499 253 529 301
rect 599 291 647 325
rect 681 291 697 325
rect 599 275 697 291
rect 745 336 775 615
rect 848 592 878 618
rect 1064 567 1094 593
rect 1187 567 1217 593
rect 1523 592 1553 618
rect 1613 592 1643 618
rect 1387 496 1417 522
rect 1064 384 1094 399
rect 1187 384 1217 399
rect 848 353 878 368
rect 1061 361 1097 384
rect 845 336 881 353
rect 745 320 881 336
rect 745 286 763 320
rect 797 286 831 320
rect 865 286 881 320
rect 599 253 629 275
rect 745 270 881 286
rect 1027 345 1131 361
rect 1027 311 1081 345
rect 1115 311 1131 345
rect 1027 295 1131 311
rect 1184 300 1220 384
rect 1387 353 1417 368
rect 1523 353 1553 368
rect 1613 353 1643 368
rect 1384 336 1420 353
rect 1339 320 1435 336
rect 1520 334 1556 353
rect 1339 300 1385 320
rect 92 55 122 81
rect 194 55 224 81
rect 299 55 329 81
rect 397 51 427 169
rect 813 237 843 270
rect 499 99 529 125
rect 599 51 629 125
rect 397 21 629 51
rect 1027 202 1057 295
rect 1190 286 1385 300
rect 1419 286 1435 320
rect 1190 270 1435 286
rect 1485 321 1558 334
rect 1610 321 1646 353
rect 1485 318 1646 321
rect 1485 284 1501 318
rect 1535 284 1646 318
rect 1190 247 1220 270
rect 1127 217 1220 247
rect 1339 246 1369 270
rect 1485 268 1646 284
rect 1528 246 1558 268
rect 1614 246 1644 268
rect 1127 202 1157 217
rect 813 63 843 89
rect 1339 136 1369 162
rect 1027 48 1057 74
rect 1127 48 1157 74
rect 1528 72 1558 98
rect 1614 72 1644 98
<< polycont >>
rect 99 263 133 297
rect 207 291 241 325
rect 647 291 681 325
rect 763 286 797 320
rect 831 286 865 320
rect 1081 311 1115 345
rect 1385 286 1419 320
rect 1501 284 1535 318
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 17 561 89 577
rect 17 527 39 561
rect 73 527 89 561
rect 17 492 89 527
rect 17 458 39 492
rect 73 458 89 492
rect 129 521 185 649
rect 129 487 132 521
rect 166 487 185 521
rect 129 461 185 487
rect 219 581 735 615
rect 219 561 275 581
rect 219 527 239 561
rect 273 527 275 561
rect 669 576 735 581
rect 17 276 65 458
rect 219 440 275 527
rect 219 424 239 440
rect 17 242 31 276
rect 99 406 239 424
rect 273 406 275 440
rect 99 390 275 406
rect 309 513 521 547
rect 669 542 685 576
rect 719 542 735 576
rect 891 597 957 649
rect 891 563 907 597
rect 941 563 957 597
rect 891 547 957 563
rect 1107 581 1442 615
rect 1107 547 1123 581
rect 1157 547 1173 581
rect 1214 531 1264 547
rect 99 297 149 390
rect 133 263 149 297
rect 191 325 263 356
rect 191 291 207 325
rect 241 291 263 325
rect 191 275 263 291
rect 309 276 343 513
rect 455 489 521 513
rect 377 441 421 479
rect 411 407 421 441
rect 377 344 421 407
rect 455 455 471 489
rect 505 455 521 489
rect 455 419 521 455
rect 455 385 471 419
rect 505 385 521 419
rect 455 378 521 385
rect 567 508 613 524
rect 1214 513 1230 531
rect 917 508 1230 513
rect 567 474 579 508
rect 613 497 1230 508
rect 613 479 1264 497
rect 613 474 951 479
rect 567 425 629 474
rect 567 391 579 425
rect 613 391 629 425
rect 567 375 629 391
rect 679 406 801 440
rect 835 406 851 440
rect 679 390 851 406
rect 377 310 551 344
rect 679 341 713 390
rect 511 276 551 310
rect 99 247 149 263
rect 17 213 65 242
rect 115 241 149 247
rect 309 242 319 276
rect 353 242 477 276
rect 17 197 81 213
rect 115 207 269 241
rect 309 239 477 242
rect 309 233 438 239
rect 17 163 47 197
rect 219 197 269 207
rect 427 205 438 233
rect 472 205 477 239
rect 17 127 81 163
rect 17 93 47 127
rect 17 77 81 93
rect 117 139 133 173
rect 167 139 183 173
rect 117 17 183 139
rect 219 163 235 197
rect 219 127 269 163
rect 219 93 235 127
rect 325 177 391 199
rect 427 187 477 205
rect 545 257 551 276
rect 631 325 713 341
rect 631 291 647 325
rect 681 291 713 325
rect 631 275 713 291
rect 545 242 597 257
rect 511 241 597 242
rect 511 207 543 241
rect 577 207 597 241
rect 511 191 597 207
rect 679 225 713 275
rect 747 320 881 356
rect 747 286 763 320
rect 797 286 831 320
rect 865 286 881 320
rect 747 270 881 286
rect 679 191 768 225
rect 802 191 818 225
rect 917 193 951 474
rect 1214 445 1264 479
rect 985 411 1017 445
rect 1051 411 1067 445
rect 985 395 1067 411
rect 1214 411 1230 445
rect 1214 395 1264 411
rect 1301 462 1374 500
rect 1301 428 1340 462
rect 985 276 1031 395
rect 1301 390 1374 428
rect 1408 424 1442 581
rect 1476 580 1510 649
rect 1476 508 1510 546
rect 1476 458 1510 474
rect 1550 580 1619 596
rect 1550 546 1566 580
rect 1600 546 1619 580
rect 1550 499 1619 546
rect 1550 465 1566 499
rect 1600 465 1619 499
rect 1408 390 1516 424
rect 1301 361 1335 390
rect 1065 345 1335 361
rect 1065 311 1081 345
rect 1115 311 1335 345
rect 1065 295 1335 311
rect 985 242 991 276
rect 1025 261 1031 276
rect 1025 242 1232 261
rect 985 227 1232 242
rect 325 143 340 177
rect 374 153 391 177
rect 917 159 982 193
rect 1016 159 1032 193
rect 917 157 1032 159
rect 511 153 1032 157
rect 374 143 1032 153
rect 325 123 1032 143
rect 325 119 545 123
rect 966 120 1032 123
rect 219 85 269 93
rect 640 85 656 89
rect 219 55 656 85
rect 690 55 706 89
rect 219 51 706 55
rect 854 55 870 89
rect 904 55 920 89
rect 966 86 982 120
rect 1016 86 1032 120
rect 966 70 1032 86
rect 1066 159 1082 193
rect 1116 159 1132 193
rect 1066 116 1132 159
rect 1166 179 1232 227
rect 1278 234 1335 295
rect 1369 320 1435 356
rect 1369 286 1385 320
rect 1419 286 1435 320
rect 1369 270 1435 286
rect 1482 334 1516 390
rect 1550 418 1619 465
rect 1550 384 1566 418
rect 1600 384 1619 418
rect 1550 368 1619 384
rect 1482 318 1551 334
rect 1482 284 1501 318
rect 1535 284 1551 318
rect 1482 268 1551 284
rect 1482 236 1516 268
rect 1278 200 1294 234
rect 1328 200 1344 234
rect 1378 202 1516 236
rect 1585 234 1619 368
rect 1656 580 1706 649
rect 1690 546 1706 580
rect 1656 497 1706 546
rect 1690 463 1706 497
rect 1656 414 1706 463
rect 1690 380 1706 414
rect 1656 364 1706 380
rect 1553 218 1619 234
rect 1166 145 1182 179
rect 1216 145 1232 179
rect 1378 166 1412 202
rect 1553 184 1569 218
rect 1603 184 1619 218
rect 1166 119 1232 145
rect 1266 132 1412 166
rect 1446 134 1462 168
rect 1496 134 1517 168
rect 1066 82 1082 116
rect 1116 85 1132 116
rect 1266 85 1300 132
rect 1446 98 1517 134
rect 1116 82 1300 85
rect 854 17 920 55
rect 1066 51 1300 82
rect 1380 82 1517 98
rect 1553 144 1619 184
rect 1553 110 1569 144
rect 1603 110 1619 144
rect 1553 88 1619 110
rect 1655 234 1705 250
rect 1689 200 1705 234
rect 1655 144 1705 200
rect 1689 110 1705 144
rect 1380 48 1396 82
rect 1430 48 1467 82
rect 1501 48 1517 82
rect 1380 17 1517 48
rect 1655 17 1705 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 242 65 276
rect 319 242 353 276
rect 511 242 545 276
rect 991 242 1025 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 19 276 77 282
rect 19 242 31 276
rect 65 273 77 276
rect 307 276 365 282
rect 307 273 319 276
rect 65 245 319 273
rect 65 242 77 245
rect 19 236 77 242
rect 307 242 319 245
rect 353 242 365 276
rect 307 236 365 242
rect 499 276 557 282
rect 499 242 511 276
rect 545 273 557 276
rect 979 276 1037 282
rect 979 273 991 276
rect 545 245 991 273
rect 545 242 557 245
rect 499 236 557 242
rect 979 242 991 245
rect 1025 242 1037 276
rect 979 236 1037 242
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xnor3_2
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 1567 94 1601 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 1567 168 1601 202 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C
port 3 nsew
flabel corelocali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1728 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 615708
string GDS_START 602552
<< end >>
