magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 737 47 767 177
rect 935 47 965 177
rect 1029 47 1059 177
rect 1123 47 1153 177
rect 1227 47 1257 177
rect 1311 47 1341 177
rect 1405 47 1435 177
rect 1499 47 1529 177
rect 1603 47 1633 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
rect 1501 297 1537 497
rect 1595 297 1631 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 95 173 177
rect 109 61 129 95
rect 163 61 173 95
rect 109 47 173 61
rect 203 163 267 177
rect 203 129 223 163
rect 257 129 267 163
rect 203 95 267 129
rect 203 61 223 95
rect 257 61 267 95
rect 203 47 267 61
rect 297 95 371 177
rect 297 61 317 95
rect 351 61 371 95
rect 297 47 371 61
rect 401 163 455 177
rect 401 129 411 163
rect 445 129 455 163
rect 401 95 455 129
rect 401 61 411 95
rect 445 61 455 95
rect 401 47 455 61
rect 485 163 549 177
rect 485 129 505 163
rect 539 129 549 163
rect 485 47 549 129
rect 579 95 643 177
rect 579 61 599 95
rect 633 61 643 95
rect 579 47 643 61
rect 673 163 737 177
rect 673 129 693 163
rect 727 129 737 163
rect 673 47 737 129
rect 767 95 829 177
rect 767 61 787 95
rect 821 61 829 95
rect 767 47 829 61
rect 883 95 935 177
rect 883 61 891 95
rect 925 61 935 95
rect 883 47 935 61
rect 965 163 1029 177
rect 965 129 985 163
rect 1019 129 1029 163
rect 965 47 1029 129
rect 1059 95 1123 177
rect 1059 61 1079 95
rect 1113 61 1123 95
rect 1059 47 1123 61
rect 1153 163 1227 177
rect 1153 129 1173 163
rect 1207 129 1227 163
rect 1153 47 1227 129
rect 1257 163 1311 177
rect 1257 129 1267 163
rect 1301 129 1311 163
rect 1257 95 1311 129
rect 1257 61 1267 95
rect 1301 61 1311 95
rect 1257 47 1311 61
rect 1341 95 1405 177
rect 1341 61 1361 95
rect 1395 61 1405 95
rect 1341 47 1405 61
rect 1435 163 1499 177
rect 1435 129 1455 163
rect 1489 129 1499 163
rect 1435 95 1499 129
rect 1435 61 1455 95
rect 1489 61 1499 95
rect 1435 47 1499 61
rect 1529 95 1603 177
rect 1529 61 1549 95
rect 1583 61 1603 95
rect 1529 47 1603 61
rect 1633 163 1685 177
rect 1633 129 1643 163
rect 1677 129 1685 163
rect 1633 95 1685 129
rect 1633 61 1643 95
rect 1677 61 1685 95
rect 1633 47 1685 61
<< pdiff >>
rect 27 481 81 497
rect 27 447 35 481
rect 69 447 81 481
rect 27 413 81 447
rect 27 379 35 413
rect 69 379 81 413
rect 27 345 81 379
rect 27 311 35 345
rect 69 311 81 345
rect 27 297 81 311
rect 117 409 175 497
rect 117 375 129 409
rect 163 375 175 409
rect 117 341 175 375
rect 117 307 129 341
rect 163 307 175 341
rect 117 297 175 307
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 297 269 375
rect 305 409 363 497
rect 305 375 317 409
rect 351 375 363 409
rect 305 341 363 375
rect 305 307 317 341
rect 351 307 363 341
rect 305 297 363 307
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 297 457 375
rect 493 409 551 497
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 477 645 497
rect 587 443 599 477
rect 633 443 645 477
rect 587 409 645 443
rect 587 375 599 409
rect 633 375 645 409
rect 587 297 645 375
rect 681 409 739 497
rect 681 375 693 409
rect 727 375 739 409
rect 681 341 739 375
rect 681 307 693 341
rect 727 307 739 341
rect 681 297 739 307
rect 775 477 937 497
rect 775 443 787 477
rect 821 443 891 477
rect 925 443 937 477
rect 775 409 937 443
rect 775 375 787 409
rect 821 375 891 409
rect 925 375 937 409
rect 775 341 937 375
rect 775 307 787 341
rect 821 307 891 341
rect 925 307 937 341
rect 775 297 937 307
rect 973 477 1031 497
rect 973 443 985 477
rect 1019 443 1031 477
rect 973 409 1031 443
rect 973 375 985 409
rect 1019 375 1031 409
rect 973 297 1031 375
rect 1067 477 1125 497
rect 1067 443 1079 477
rect 1113 443 1125 477
rect 1067 409 1125 443
rect 1067 375 1079 409
rect 1113 375 1125 409
rect 1067 341 1125 375
rect 1067 307 1079 341
rect 1113 307 1125 341
rect 1067 297 1125 307
rect 1161 477 1219 497
rect 1161 443 1173 477
rect 1207 443 1219 477
rect 1161 409 1219 443
rect 1161 375 1173 409
rect 1207 375 1219 409
rect 1161 297 1219 375
rect 1255 477 1313 497
rect 1255 443 1267 477
rect 1301 443 1313 477
rect 1255 409 1313 443
rect 1255 375 1267 409
rect 1301 375 1313 409
rect 1255 341 1313 375
rect 1255 307 1267 341
rect 1301 307 1313 341
rect 1255 297 1313 307
rect 1349 477 1407 497
rect 1349 443 1361 477
rect 1395 443 1407 477
rect 1349 409 1407 443
rect 1349 375 1361 409
rect 1395 375 1407 409
rect 1349 297 1407 375
rect 1443 477 1501 497
rect 1443 443 1455 477
rect 1489 443 1501 477
rect 1443 409 1501 443
rect 1443 375 1455 409
rect 1489 375 1501 409
rect 1443 341 1501 375
rect 1443 307 1455 341
rect 1489 307 1501 341
rect 1443 297 1501 307
rect 1537 477 1595 497
rect 1537 443 1549 477
rect 1583 443 1595 477
rect 1537 409 1595 443
rect 1537 375 1549 409
rect 1583 375 1595 409
rect 1537 297 1595 375
rect 1631 477 1693 497
rect 1631 443 1643 477
rect 1677 443 1693 477
rect 1631 409 1693 443
rect 1631 375 1643 409
rect 1677 375 1693 409
rect 1631 341 1693 375
rect 1631 307 1643 341
rect 1677 307 1693 341
rect 1631 297 1693 307
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 61 163 95
rect 223 129 257 163
rect 223 61 257 95
rect 317 61 351 95
rect 411 129 445 163
rect 411 61 445 95
rect 505 129 539 163
rect 599 61 633 95
rect 693 129 727 163
rect 787 61 821 95
rect 891 61 925 95
rect 985 129 1019 163
rect 1079 61 1113 95
rect 1173 129 1207 163
rect 1267 129 1301 163
rect 1267 61 1301 95
rect 1361 61 1395 95
rect 1455 129 1489 163
rect 1455 61 1489 95
rect 1549 61 1583 95
rect 1643 129 1677 163
rect 1643 61 1677 95
<< pdiffc >>
rect 35 447 69 481
rect 35 379 69 413
rect 35 311 69 345
rect 129 375 163 409
rect 129 307 163 341
rect 223 443 257 477
rect 223 375 257 409
rect 317 375 351 409
rect 317 307 351 341
rect 411 443 445 477
rect 411 375 445 409
rect 505 375 539 409
rect 505 307 539 341
rect 599 443 633 477
rect 599 375 633 409
rect 693 375 727 409
rect 693 307 727 341
rect 787 443 821 477
rect 891 443 925 477
rect 787 375 821 409
rect 891 375 925 409
rect 787 307 821 341
rect 891 307 925 341
rect 985 443 1019 477
rect 985 375 1019 409
rect 1079 443 1113 477
rect 1079 375 1113 409
rect 1079 307 1113 341
rect 1173 443 1207 477
rect 1173 375 1207 409
rect 1267 443 1301 477
rect 1267 375 1301 409
rect 1267 307 1301 341
rect 1361 443 1395 477
rect 1361 375 1395 409
rect 1455 443 1489 477
rect 1455 375 1489 409
rect 1455 307 1489 341
rect 1549 443 1583 477
rect 1549 375 1583 409
rect 1643 443 1677 477
rect 1643 375 1677 409
rect 1643 307 1677 341
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 1501 497 1537 523
rect 1595 497 1631 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 1501 282 1537 297
rect 1595 282 1631 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 79 249 401 265
rect 79 215 107 249
rect 141 215 185 249
rect 219 215 263 249
rect 297 215 341 249
rect 375 215 401 249
rect 79 199 401 215
rect 79 177 109 199
rect 173 177 203 199
rect 267 177 297 199
rect 371 177 401 199
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 935 265 975 282
rect 1029 265 1069 282
rect 1123 265 1163 282
rect 1217 265 1257 282
rect 455 249 812 265
rect 455 215 606 249
rect 640 215 684 249
rect 718 215 752 249
rect 786 215 812 249
rect 455 199 812 215
rect 935 249 1257 265
rect 935 215 951 249
rect 985 215 1029 249
rect 1063 215 1107 249
rect 1141 215 1185 249
rect 1219 215 1257 249
rect 935 199 1257 215
rect 455 177 485 199
rect 549 177 579 199
rect 643 177 673 199
rect 737 177 767 199
rect 935 177 965 199
rect 1029 177 1059 199
rect 1123 177 1153 199
rect 1227 177 1257 199
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 1499 265 1539 282
rect 1593 265 1633 282
rect 1311 249 1633 265
rect 1311 215 1327 249
rect 1361 215 1405 249
rect 1439 215 1483 249
rect 1517 215 1561 249
rect 1595 215 1633 249
rect 1311 199 1633 215
rect 1311 177 1341 199
rect 1405 177 1435 199
rect 1499 177 1529 199
rect 1603 177 1633 199
rect 79 21 109 47
rect 173 21 203 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 737 21 767 47
rect 935 21 965 47
rect 1029 21 1059 47
rect 1123 21 1153 47
rect 1227 21 1257 47
rect 1311 21 1341 47
rect 1405 21 1435 47
rect 1499 21 1529 47
rect 1603 21 1633 47
<< polycont >>
rect 107 215 141 249
rect 185 215 219 249
rect 263 215 297 249
rect 341 215 375 249
rect 606 215 640 249
rect 684 215 718 249
rect 752 215 786 249
rect 951 215 985 249
rect 1029 215 1063 249
rect 1107 215 1141 249
rect 1185 215 1219 249
rect 1327 215 1361 249
rect 1405 215 1439 249
rect 1483 215 1517 249
rect 1561 215 1595 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 481 933 493
rect 18 447 35 481
rect 69 477 933 481
rect 69 459 223 477
rect 69 447 85 459
rect 18 413 85 447
rect 215 443 223 459
rect 257 459 411 477
rect 257 443 265 459
rect 18 379 35 413
rect 69 379 85 413
rect 18 345 85 379
rect 18 311 35 345
rect 69 311 85 345
rect 18 291 85 311
rect 129 409 171 425
rect 163 375 171 409
rect 129 341 171 375
rect 215 409 265 443
rect 403 443 411 459
rect 445 459 599 477
rect 445 443 453 459
rect 215 375 223 409
rect 257 375 265 409
rect 215 359 265 375
rect 309 409 359 425
rect 309 375 317 409
rect 351 375 359 409
rect 163 325 171 341
rect 309 341 359 375
rect 403 409 453 443
rect 591 443 599 459
rect 633 459 787 477
rect 633 443 641 459
rect 403 375 411 409
rect 445 375 453 409
rect 403 359 453 375
rect 497 409 547 425
rect 497 375 505 409
rect 539 375 547 409
rect 309 325 317 341
rect 163 307 317 325
rect 351 325 359 341
rect 497 341 547 375
rect 591 409 641 443
rect 779 443 787 459
rect 821 443 891 477
rect 925 443 933 477
rect 591 375 599 409
rect 633 375 641 409
rect 591 359 641 375
rect 685 409 735 425
rect 685 375 693 409
rect 727 375 735 409
rect 497 325 505 341
rect 351 307 505 325
rect 539 325 547 341
rect 685 341 735 375
rect 685 325 693 341
rect 539 307 693 325
rect 727 307 735 341
rect 129 289 735 307
rect 779 409 933 443
rect 779 375 787 409
rect 821 375 891 409
rect 925 375 933 409
rect 779 341 933 375
rect 977 477 1027 527
rect 977 443 985 477
rect 1019 443 1027 477
rect 977 409 1027 443
rect 977 375 985 409
rect 1019 375 1027 409
rect 977 359 1027 375
rect 1071 477 1121 493
rect 1071 443 1079 477
rect 1113 443 1121 477
rect 1071 409 1121 443
rect 1071 375 1079 409
rect 1113 375 1121 409
rect 779 307 787 341
rect 821 307 891 341
rect 925 325 933 341
rect 1071 341 1121 375
rect 1165 477 1215 527
rect 1165 443 1173 477
rect 1207 443 1215 477
rect 1165 409 1215 443
rect 1165 375 1173 409
rect 1207 375 1215 409
rect 1165 359 1215 375
rect 1259 477 1309 493
rect 1259 443 1267 477
rect 1301 443 1309 477
rect 1259 409 1309 443
rect 1259 375 1267 409
rect 1301 375 1309 409
rect 1071 325 1079 341
rect 925 307 1079 325
rect 1113 325 1121 341
rect 1259 341 1309 375
rect 1353 477 1403 527
rect 1353 443 1361 477
rect 1395 443 1403 477
rect 1353 409 1403 443
rect 1353 375 1361 409
rect 1395 375 1403 409
rect 1353 359 1403 375
rect 1447 477 1497 493
rect 1447 443 1455 477
rect 1489 443 1497 477
rect 1447 409 1497 443
rect 1447 375 1455 409
rect 1489 375 1497 409
rect 1259 325 1267 341
rect 1113 307 1267 325
rect 1301 325 1309 341
rect 1447 341 1497 375
rect 1541 477 1591 527
rect 1541 443 1549 477
rect 1583 443 1591 477
rect 1541 409 1591 443
rect 1541 375 1549 409
rect 1583 375 1591 409
rect 1541 359 1591 375
rect 1635 477 1685 493
rect 1635 443 1643 477
rect 1677 443 1685 477
rect 1635 409 1685 443
rect 1635 375 1643 409
rect 1677 375 1685 409
rect 1447 325 1455 341
rect 1301 307 1455 325
rect 1489 325 1497 341
rect 1635 341 1685 375
rect 1635 325 1643 341
rect 1489 307 1643 325
rect 1677 307 1685 341
rect 779 291 1685 307
rect 18 249 419 255
rect 18 215 107 249
rect 141 215 185 249
rect 219 215 263 249
rect 297 215 341 249
rect 375 215 419 249
rect 19 163 445 181
rect 19 129 35 163
rect 69 145 223 163
rect 69 129 85 145
rect 19 95 85 129
rect 197 129 223 145
rect 257 145 411 163
rect 257 129 273 145
rect 19 61 35 95
rect 69 61 85 95
rect 19 51 85 61
rect 129 95 163 111
rect 129 17 163 61
rect 197 95 273 129
rect 385 129 411 145
rect 479 177 539 289
rect 573 249 888 255
rect 573 215 606 249
rect 640 215 684 249
rect 718 215 752 249
rect 786 215 888 249
rect 935 249 1257 257
rect 935 215 951 249
rect 985 215 1029 249
rect 1063 215 1107 249
rect 1141 215 1185 249
rect 1219 215 1257 249
rect 1302 249 1707 257
rect 1302 215 1327 249
rect 1361 215 1405 249
rect 1439 215 1483 249
rect 1517 215 1561 249
rect 1595 215 1707 249
rect 479 163 1223 177
rect 479 129 505 163
rect 539 129 693 163
rect 727 129 985 163
rect 1019 129 1173 163
rect 1207 129 1223 163
rect 1267 163 1693 181
rect 1301 145 1455 163
rect 1301 129 1317 145
rect 197 61 223 95
rect 257 61 273 95
rect 197 51 273 61
rect 317 95 351 111
rect 317 17 351 61
rect 385 95 445 129
rect 1267 95 1317 129
rect 1429 129 1455 145
rect 1489 145 1643 163
rect 1489 129 1505 145
rect 385 61 411 95
rect 445 61 599 95
rect 633 61 787 95
rect 821 61 837 95
rect 385 51 837 61
rect 875 61 891 95
rect 925 61 1079 95
rect 1113 61 1267 95
rect 1301 61 1317 95
rect 875 51 1317 61
rect 1361 95 1395 111
rect 1361 17 1395 61
rect 1429 95 1505 129
rect 1617 129 1643 145
rect 1677 129 1693 163
rect 1429 61 1455 95
rect 1489 61 1505 95
rect 1429 51 1505 61
rect 1549 95 1583 111
rect 1549 17 1583 61
rect 1617 95 1693 129
rect 1617 61 1643 95
rect 1677 61 1693 95
rect 1617 51 1693 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel corelocali s 1339 238 1339 238 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel corelocali s 217 221 251 255 0 FreeSans 400 180 0 0 B2
port 4 nsew
flabel corelocali s 971 238 971 238 0 FreeSans 400 0 0 0 A1
port 1 nsew
flabel corelocali s 599 238 599 238 0 FreeSans 400 180 0 0 B1
port 3 nsew
flabel corelocali s 132 289 166 323 0 FreeSans 400 180 0 0 Y
port 9 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1304530
string GDS_START 1291812
<< end >>
