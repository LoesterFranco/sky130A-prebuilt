magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 17 165 69 490
rect 187 199 257 323
rect 295 199 387 323
rect 435 199 531 323
rect 565 199 645 323
rect 17 131 415 165
rect 181 60 221 131
rect 375 62 415 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 465 437 541 527
rect 105 359 713 401
rect 105 199 149 359
rect 679 165 713 359
rect 71 17 137 96
rect 265 17 331 97
rect 449 17 547 165
rect 618 131 713 165
rect 618 81 652 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 435 199 531 323 6 A
port 1 nsew signal input
rlabel locali s 295 199 387 323 6 B
port 2 nsew signal input
rlabel locali s 187 199 257 323 6 C
port 3 nsew signal input
rlabel locali s 565 199 645 323 6 D_N
port 4 nsew signal input
rlabel locali s 375 62 415 131 6 Y
port 5 nsew signal output
rlabel locali s 181 60 221 131 6 Y
port 5 nsew signal output
rlabel locali s 17 165 69 490 6 Y
port 5 nsew signal output
rlabel locali s 17 131 415 165 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2506440
string GDS_START 2500946
<< end >>
