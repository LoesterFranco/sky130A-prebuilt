magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 202 394 268 596
rect 382 394 448 596
rect 133 360 448 394
rect 133 356 167 360
rect 25 226 167 356
rect 511 270 570 356
rect 25 192 409 226
rect 672 270 737 356
rect 1081 252 1223 356
rect 1273 252 1415 356
rect 187 70 237 192
rect 359 70 409 192
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 112 428 162 649
rect 308 428 342 649
rect 482 390 556 649
rect 658 424 724 596
rect 812 581 1042 615
rect 812 458 878 581
rect 604 390 830 424
rect 207 260 477 326
rect 443 236 477 260
rect 443 202 563 236
rect 604 226 638 390
rect 771 294 830 390
rect 913 236 952 547
rect 992 424 1042 581
rect 1082 458 1132 649
rect 1172 424 1238 596
rect 1278 458 1312 649
rect 1352 424 1418 596
rect 992 390 1418 424
rect 101 17 151 158
rect 273 17 323 158
rect 445 17 495 168
rect 529 85 563 202
rect 597 119 638 226
rect 672 202 963 236
rect 672 85 706 202
rect 529 51 706 85
rect 740 17 877 168
rect 913 120 963 202
rect 1001 184 1419 218
rect 1001 154 1223 184
rect 913 70 1153 120
rect 1189 70 1223 154
rect 1259 70 1333 150
rect 1369 70 1419 184
rect 1299 17 1333 70
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel locali s 511 270 570 356 6 A1_N
port 1 nsew signal input
rlabel locali s 672 270 737 356 6 A2_N
port 2 nsew signal input
rlabel locali s 1273 252 1415 356 6 B1
port 3 nsew signal input
rlabel locali s 1081 252 1223 356 6 B2
port 4 nsew signal input
rlabel locali s 382 394 448 596 6 X
port 5 nsew signal output
rlabel locali s 359 70 409 192 6 X
port 5 nsew signal output
rlabel locali s 202 394 268 596 6 X
port 5 nsew signal output
rlabel locali s 187 70 237 192 6 X
port 5 nsew signal output
rlabel locali s 133 360 448 394 6 X
port 5 nsew signal output
rlabel locali s 133 356 167 360 6 X
port 5 nsew signal output
rlabel locali s 25 226 167 356 6 X
port 5 nsew signal output
rlabel locali s 25 192 409 226 6 X
port 5 nsew signal output
rlabel metal1 s 0 -49 1440 49 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1440 715 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3651272
string GDS_START 3639722
<< end >>
