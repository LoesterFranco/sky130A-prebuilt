magic
tech sky130A
magscale 1 2
timestamp 1599588205
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 287 47 317 177
rect 381 47 411 177
rect 475 47 505 177
rect 569 47 599 177
rect 653 47 683 177
rect 747 47 777 177
rect 841 47 871 177
rect 945 47 975 177
rect 1143 47 1173 177
rect 1237 47 1267 177
rect 1331 47 1361 177
rect 1425 47 1455 177
<< pmoshvt >>
rect 81 297 117 497
rect 279 297 315 497
rect 373 297 409 497
rect 467 297 503 497
rect 561 297 597 497
rect 655 297 691 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1135 297 1171 497
rect 1229 297 1265 497
rect 1323 297 1359 497
rect 1417 297 1453 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 171 177
rect 109 59 129 93
rect 163 59 171 93
rect 109 47 171 59
rect 225 93 287 177
rect 225 59 233 93
rect 267 59 287 93
rect 225 47 287 59
rect 317 161 381 177
rect 317 127 327 161
rect 361 127 381 161
rect 317 47 381 127
rect 411 93 475 177
rect 411 59 421 93
rect 455 59 475 93
rect 411 47 475 59
rect 505 161 569 177
rect 505 127 515 161
rect 549 127 569 161
rect 505 47 569 127
rect 599 93 653 177
rect 599 59 609 93
rect 643 59 653 93
rect 599 47 653 59
rect 683 161 747 177
rect 683 127 703 161
rect 737 127 747 161
rect 683 47 747 127
rect 777 93 841 177
rect 777 59 797 93
rect 831 59 841 93
rect 777 47 841 59
rect 871 161 945 177
rect 871 127 891 161
rect 925 127 945 161
rect 871 47 945 127
rect 975 93 1027 177
rect 975 59 985 93
rect 1019 59 1027 93
rect 975 47 1027 59
rect 1081 93 1143 177
rect 1081 59 1089 93
rect 1123 59 1143 93
rect 1081 47 1143 59
rect 1173 161 1237 177
rect 1173 127 1183 161
rect 1217 127 1237 161
rect 1173 93 1237 127
rect 1173 59 1183 93
rect 1217 59 1237 93
rect 1173 47 1237 59
rect 1267 93 1331 177
rect 1267 59 1277 93
rect 1311 59 1331 93
rect 1267 47 1331 59
rect 1361 161 1425 177
rect 1361 127 1371 161
rect 1405 127 1425 161
rect 1361 93 1425 127
rect 1361 59 1371 93
rect 1405 59 1425 93
rect 1361 47 1425 59
rect 1455 161 1527 177
rect 1455 127 1481 161
rect 1515 127 1527 161
rect 1455 93 1527 127
rect 1455 59 1481 93
rect 1515 59 1527 93
rect 1455 47 1527 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 171 497
rect 117 451 129 485
rect 163 451 171 485
rect 117 417 171 451
rect 117 383 129 417
rect 163 383 171 417
rect 117 349 171 383
rect 117 315 129 349
rect 163 315 171 349
rect 117 297 171 315
rect 225 485 279 497
rect 225 451 233 485
rect 267 451 279 485
rect 225 417 279 451
rect 225 383 233 417
rect 267 383 279 417
rect 225 349 279 383
rect 225 315 233 349
rect 267 315 279 349
rect 225 297 279 315
rect 315 485 373 497
rect 315 451 327 485
rect 361 451 373 485
rect 315 417 373 451
rect 315 383 327 417
rect 361 383 373 417
rect 315 349 373 383
rect 315 315 327 349
rect 361 315 373 349
rect 315 297 373 315
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 297 467 383
rect 503 485 561 497
rect 503 451 515 485
rect 549 451 561 485
rect 503 417 561 451
rect 503 383 515 417
rect 549 383 561 417
rect 503 349 561 383
rect 503 315 515 349
rect 549 315 561 349
rect 503 297 561 315
rect 597 485 655 497
rect 597 451 609 485
rect 643 451 655 485
rect 597 297 655 451
rect 691 485 749 497
rect 691 451 703 485
rect 737 451 749 485
rect 691 417 749 451
rect 691 383 703 417
rect 737 383 749 417
rect 691 349 749 383
rect 691 315 703 349
rect 737 315 749 349
rect 691 297 749 315
rect 785 485 843 497
rect 785 451 797 485
rect 831 451 843 485
rect 785 417 843 451
rect 785 383 797 417
rect 831 383 843 417
rect 785 297 843 383
rect 879 485 937 497
rect 879 451 891 485
rect 925 451 937 485
rect 879 417 937 451
rect 879 383 891 417
rect 925 383 937 417
rect 879 349 937 383
rect 879 315 891 349
rect 925 315 937 349
rect 879 297 937 315
rect 973 485 1027 497
rect 973 451 985 485
rect 1019 451 1027 485
rect 973 417 1027 451
rect 973 383 985 417
rect 1019 383 1027 417
rect 973 297 1027 383
rect 1081 485 1135 497
rect 1081 451 1089 485
rect 1123 451 1135 485
rect 1081 417 1135 451
rect 1081 383 1089 417
rect 1123 383 1135 417
rect 1081 297 1135 383
rect 1171 485 1229 497
rect 1171 451 1183 485
rect 1217 451 1229 485
rect 1171 417 1229 451
rect 1171 383 1183 417
rect 1217 383 1229 417
rect 1171 349 1229 383
rect 1171 315 1183 349
rect 1217 315 1229 349
rect 1171 297 1229 315
rect 1265 485 1323 497
rect 1265 451 1277 485
rect 1311 451 1323 485
rect 1265 417 1323 451
rect 1265 383 1277 417
rect 1311 383 1323 417
rect 1265 297 1323 383
rect 1359 485 1417 497
rect 1359 451 1371 485
rect 1405 451 1417 485
rect 1359 417 1417 451
rect 1359 383 1371 417
rect 1405 383 1417 417
rect 1359 349 1417 383
rect 1359 315 1371 349
rect 1405 315 1417 349
rect 1359 297 1417 315
rect 1453 485 1527 497
rect 1453 451 1481 485
rect 1515 451 1527 485
rect 1453 417 1527 451
rect 1453 383 1481 417
rect 1515 383 1527 417
rect 1453 349 1527 383
rect 1453 315 1481 349
rect 1515 315 1527 349
rect 1453 297 1527 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 233 59 267 93
rect 327 127 361 161
rect 421 59 455 93
rect 515 127 549 161
rect 609 59 643 93
rect 703 127 737 161
rect 797 59 831 93
rect 891 127 925 161
rect 985 59 1019 93
rect 1089 59 1123 93
rect 1183 127 1217 161
rect 1183 59 1217 93
rect 1277 59 1311 93
rect 1371 127 1405 161
rect 1371 59 1405 93
rect 1481 127 1515 161
rect 1481 59 1515 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 233 451 267 485
rect 233 383 267 417
rect 233 315 267 349
rect 327 451 361 485
rect 327 383 361 417
rect 327 315 361 349
rect 421 451 455 485
rect 421 383 455 417
rect 515 451 549 485
rect 515 383 549 417
rect 515 315 549 349
rect 609 451 643 485
rect 703 451 737 485
rect 703 383 737 417
rect 703 315 737 349
rect 797 451 831 485
rect 797 383 831 417
rect 891 451 925 485
rect 891 383 925 417
rect 891 315 925 349
rect 985 451 1019 485
rect 985 383 1019 417
rect 1089 451 1123 485
rect 1089 383 1123 417
rect 1183 451 1217 485
rect 1183 383 1217 417
rect 1183 315 1217 349
rect 1277 451 1311 485
rect 1277 383 1311 417
rect 1371 451 1405 485
rect 1371 383 1405 417
rect 1371 315 1405 349
rect 1481 451 1515 485
rect 1481 383 1515 417
rect 1481 315 1515 349
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 373 497 409 523
rect 467 497 503 523
rect 561 497 597 523
rect 655 497 691 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1135 497 1171 523
rect 1229 497 1265 523
rect 1323 497 1359 523
rect 1417 497 1453 523
rect 81 282 117 297
rect 279 282 315 297
rect 373 282 409 297
rect 467 282 503 297
rect 561 282 597 297
rect 655 282 691 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1135 282 1171 297
rect 1229 282 1265 297
rect 1323 282 1359 297
rect 1417 282 1453 297
rect 79 261 119 282
rect 79 249 162 261
rect 277 259 317 282
rect 371 259 411 282
rect 465 259 505 282
rect 559 259 599 282
rect 79 215 102 249
rect 136 215 162 249
rect 79 203 162 215
rect 211 249 599 259
rect 211 215 227 249
rect 261 215 327 249
rect 361 215 421 249
rect 455 215 515 249
rect 549 215 599 249
rect 211 205 599 215
rect 79 177 109 203
rect 287 177 317 205
rect 381 177 411 205
rect 475 177 505 205
rect 569 177 599 205
rect 653 259 693 282
rect 747 259 787 282
rect 841 259 881 282
rect 935 259 975 282
rect 1133 259 1173 282
rect 1227 259 1267 282
rect 1321 259 1361 282
rect 1415 259 1455 282
rect 653 249 975 259
rect 653 215 765 249
rect 799 215 886 249
rect 920 215 975 249
rect 653 205 975 215
rect 1067 249 1455 259
rect 1067 215 1083 249
rect 1117 215 1183 249
rect 1217 215 1277 249
rect 1311 215 1370 249
rect 1404 215 1455 249
rect 1067 205 1455 215
rect 653 177 683 205
rect 747 177 777 205
rect 841 177 871 205
rect 945 177 975 205
rect 1143 177 1173 205
rect 1237 177 1267 205
rect 1331 177 1361 205
rect 1425 177 1455 205
rect 79 21 109 47
rect 287 21 317 47
rect 381 21 411 47
rect 475 21 505 47
rect 569 21 599 47
rect 653 21 683 47
rect 747 21 777 47
rect 841 21 871 47
rect 945 21 975 47
rect 1143 21 1173 47
rect 1237 21 1267 47
rect 1331 21 1361 47
rect 1425 21 1455 47
<< polycont >>
rect 102 215 136 249
rect 227 215 261 249
rect 327 215 361 249
rect 421 215 455 249
rect 515 215 549 249
rect 765 215 799 249
rect 886 215 920 249
rect 1083 215 1117 249
rect 1183 215 1217 249
rect 1277 215 1311 249
rect 1370 215 1404 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 485 85 493
rect 17 451 35 485
rect 69 451 85 485
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 17 315 35 349
rect 69 315 85 349
rect 17 289 85 315
rect 129 485 267 527
rect 163 451 233 485
rect 129 417 267 451
rect 163 383 233 417
rect 129 349 267 383
rect 163 315 233 349
rect 129 289 267 315
rect 301 485 377 493
rect 301 451 327 485
rect 361 451 377 485
rect 301 417 377 451
rect 301 383 327 417
rect 361 383 377 417
rect 301 349 377 383
rect 421 485 455 527
rect 421 417 455 451
rect 421 367 455 383
rect 489 485 565 493
rect 489 451 515 485
rect 549 451 565 485
rect 489 417 565 451
rect 609 485 643 527
rect 609 435 643 451
rect 677 485 753 493
rect 677 451 703 485
rect 737 451 753 485
rect 489 383 515 417
rect 549 401 565 417
rect 677 417 753 451
rect 677 401 703 417
rect 549 383 703 401
rect 737 383 753 417
rect 301 315 327 349
rect 361 333 377 349
rect 489 349 753 383
rect 797 485 831 527
rect 797 417 831 451
rect 797 367 831 383
rect 865 485 941 493
rect 865 451 891 485
rect 925 451 941 485
rect 865 417 941 451
rect 865 383 891 417
rect 925 383 941 417
rect 489 333 515 349
rect 361 315 515 333
rect 549 315 703 349
rect 737 333 753 349
rect 865 349 941 383
rect 985 485 1123 527
rect 1019 451 1089 485
rect 985 417 1123 451
rect 1019 383 1089 417
rect 985 367 1123 383
rect 1157 485 1233 493
rect 1157 451 1183 485
rect 1217 451 1233 485
rect 1157 417 1233 451
rect 1157 383 1183 417
rect 1217 383 1233 417
rect 865 333 891 349
rect 737 315 891 333
rect 925 333 941 349
rect 1157 349 1233 383
rect 1277 485 1311 527
rect 1277 417 1311 451
rect 1277 367 1311 383
rect 1345 485 1421 493
rect 1345 451 1371 485
rect 1405 451 1421 485
rect 1345 417 1421 451
rect 1345 383 1371 417
rect 1405 383 1421 417
rect 1157 333 1183 349
rect 925 315 1183 333
rect 1217 333 1233 349
rect 1345 349 1421 383
rect 1345 333 1371 349
rect 1217 315 1371 333
rect 1405 315 1421 349
rect 301 289 1421 315
rect 1465 485 1531 527
rect 1465 451 1481 485
rect 1515 451 1531 485
rect 1465 417 1531 451
rect 1465 383 1481 417
rect 1515 383 1531 417
rect 1465 349 1531 383
rect 1465 315 1481 349
rect 1515 315 1531 349
rect 1465 289 1531 315
rect 17 181 52 289
rect 86 249 166 255
rect 86 215 102 249
rect 136 215 166 249
rect 211 249 565 255
rect 211 215 227 249
rect 261 215 327 249
rect 361 215 421 249
rect 455 215 515 249
rect 549 215 565 249
rect 609 215 711 289
rect 745 249 986 255
rect 745 215 765 249
rect 799 215 886 249
rect 920 215 986 249
rect 1037 249 1420 255
rect 1037 215 1083 249
rect 1117 215 1183 249
rect 1217 215 1277 249
rect 1311 215 1370 249
rect 1404 215 1420 249
rect 211 181 267 215
rect 609 181 643 215
rect 17 161 267 181
rect 17 127 35 161
rect 69 143 267 161
rect 301 161 643 181
rect 69 127 85 143
rect 301 127 327 161
rect 361 127 515 161
rect 549 127 643 161
rect 677 161 1421 181
rect 677 127 703 161
rect 737 127 891 161
rect 925 143 1183 161
rect 925 127 1035 143
rect 1157 127 1183 143
rect 1217 143 1371 161
rect 1217 127 1233 143
rect 17 93 85 127
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 129 93 179 109
rect 1073 93 1123 109
rect 163 59 179 93
rect 129 17 179 59
rect 217 59 233 93
rect 267 59 421 93
rect 455 59 609 93
rect 643 59 797 93
rect 831 59 985 93
rect 1019 59 1035 93
rect 217 51 1035 59
rect 1073 59 1089 93
rect 1073 17 1123 59
rect 1157 93 1233 127
rect 1345 127 1371 143
rect 1405 127 1421 161
rect 1157 59 1183 93
rect 1217 59 1233 93
rect 1157 51 1233 59
rect 1277 93 1311 109
rect 1277 17 1311 59
rect 1345 93 1421 127
rect 1345 59 1371 93
rect 1405 59 1421 93
rect 1345 51 1421 59
rect 1465 161 1531 181
rect 1465 127 1481 161
rect 1515 127 1531 161
rect 1465 93 1531 127
rect 1465 59 1481 93
rect 1515 59 1531 93
rect 1465 17 1531 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel corelocali s 121 221 155 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel corelocali s 673 221 707 255 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 949 221 983 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 765 221 799 255 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel corelocali s 673 357 707 391 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 1317 221 1351 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 1041 221 1075 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 1133 221 1167 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 1225 221 1259 255 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel corelocali s 673 289 707 323 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 nand3b_4
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2287458
string GDS_START 2275096
<< end >>
