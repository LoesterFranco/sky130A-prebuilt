magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 119 367 185 527
rect 17 211 112 265
rect 528 352 608 527
rect 642 352 719 493
rect 119 17 182 109
rect 673 109 719 352
rect 542 17 608 109
rect 642 57 719 109
rect 0 -17 736 17
<< obsli1 >>
rect 17 333 85 493
rect 277 367 352 493
rect 17 299 243 333
rect 146 177 243 299
rect 17 143 243 177
rect 318 250 352 367
rect 386 318 482 493
rect 386 284 639 318
rect 318 211 537 250
rect 318 165 352 211
rect 571 177 639 284
rect 17 51 85 143
rect 277 51 352 165
rect 386 143 639 177
rect 386 51 452 143
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 17 211 112 265 6 A
port 1 nsew signal input
rlabel locali s 673 109 719 352 6 X
port 2 nsew signal output
rlabel locali s 642 352 719 493 6 X
port 2 nsew signal output
rlabel locali s 642 57 719 109 6 X
port 2 nsew signal output
rlabel locali s 542 17 608 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 119 17 182 109 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 528 352 608 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 119 367 185 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3155080
string GDS_START 3148960
<< end >>
