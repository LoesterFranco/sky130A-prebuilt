magic
tech sky130A
magscale 1 2
timestamp 1599588238
<< locali >>
rect 23 458 89 596
rect 23 226 57 458
rect 217 290 316 356
rect 23 70 75 226
rect 374 238 455 356
rect 494 244 560 578
rect 601 260 674 578
rect 722 270 839 430
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 123 458 308 649
rect 350 424 416 569
rect 91 390 416 424
rect 91 270 157 390
rect 123 256 157 270
rect 123 222 301 256
rect 752 464 841 649
rect 109 17 189 188
rect 235 70 301 222
rect 775 204 841 206
rect 335 170 841 204
rect 335 70 401 170
rect 435 17 501 136
rect 535 70 601 170
rect 635 17 741 136
rect 775 70 841 170
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 722 270 839 430 6 A1
port 1 nsew signal input
rlabel locali s 601 260 674 578 6 A2
port 2 nsew signal input
rlabel locali s 494 244 560 578 6 A3
port 3 nsew signal input
rlabel locali s 374 238 455 356 6 A4
port 4 nsew signal input
rlabel locali s 217 290 316 356 6 B1
port 5 nsew signal input
rlabel locali s 23 458 89 596 6 X
port 6 nsew signal output
rlabel locali s 23 226 57 458 6 X
port 6 nsew signal output
rlabel locali s 23 70 75 226 6 X
port 6 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 617 864 715 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 901408
string GDS_START 893136
<< end >>
