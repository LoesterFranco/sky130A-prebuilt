magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 25 200 99 434
rect 409 346 455 356
rect 359 264 455 346
rect 2130 70 2196 596
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 21 504 87 649
rect 127 526 167 596
rect 203 546 269 649
rect 391 548 457 649
rect 127 521 174 526
rect 609 523 665 545
rect 481 521 665 523
rect 127 512 178 521
rect 478 519 665 521
rect 475 518 665 519
rect 473 517 665 518
rect 471 516 665 517
rect 469 515 665 516
rect 466 514 665 515
rect 281 512 665 514
rect 127 504 665 512
rect 699 514 850 550
rect 884 548 950 649
rect 699 505 1057 514
rect 133 489 665 504
rect 133 488 497 489
rect 133 487 494 488
rect 133 486 492 487
rect 133 484 488 486
rect 133 481 484 484
rect 133 479 481 481
rect 589 480 665 489
rect 787 480 1057 505
rect 133 476 477 479
rect 133 471 472 476
rect 589 475 674 480
rect 622 471 674 475
rect 133 466 468 471
rect 133 166 167 466
rect 506 446 555 455
rect 622 446 753 471
rect 503 441 555 446
rect 201 424 257 430
rect 201 390 223 424
rect 201 228 257 390
rect 291 380 373 432
rect 503 416 588 441
rect 640 437 753 446
rect 503 407 602 416
rect 503 397 619 407
rect 503 389 685 397
rect 562 380 685 389
rect 291 230 325 380
rect 503 310 537 355
rect 489 230 537 310
rect 291 195 537 230
rect 573 325 685 380
rect 291 194 508 195
rect 26 132 167 166
rect 26 74 92 132
rect 201 17 257 166
rect 291 70 375 194
rect 573 161 614 325
rect 719 278 753 437
rect 664 244 753 278
rect 664 209 698 244
rect 787 210 821 480
rect 923 464 1057 480
rect 419 17 485 160
rect 519 100 614 161
rect 648 134 698 209
rect 732 134 821 210
rect 855 225 889 425
rect 923 315 957 464
rect 991 424 1057 430
rect 1025 390 1057 424
rect 991 359 1057 390
rect 1103 349 1169 649
rect 1203 371 1269 551
rect 1303 495 1525 561
rect 923 259 1137 315
rect 1203 226 1237 371
rect 1303 337 1337 495
rect 1171 225 1237 226
rect 855 191 1237 225
rect 861 123 1137 157
rect 861 100 895 123
rect 519 66 895 100
rect 984 17 1069 89
rect 1103 85 1137 123
rect 1171 119 1237 191
rect 1271 303 1337 337
rect 1271 169 1305 303
rect 1391 269 1457 461
rect 1491 346 1525 495
rect 1559 489 1625 649
rect 1659 489 1777 555
rect 1818 489 1884 649
rect 1743 455 1777 489
rect 1561 424 1679 455
rect 1561 390 1567 424
rect 1601 390 1679 424
rect 1743 421 1875 455
rect 1561 384 1679 390
rect 1741 346 1807 378
rect 1491 312 1807 346
rect 1841 278 1875 421
rect 1918 406 1984 581
rect 1345 203 1491 269
rect 1525 244 1875 278
rect 1932 326 1984 406
rect 2030 364 2096 649
rect 1932 260 2038 326
rect 1525 212 1591 244
rect 1271 119 1423 169
rect 1457 85 1491 203
rect 1103 51 1491 85
rect 1554 17 1638 143
rect 1736 77 1802 244
rect 1846 17 1896 210
rect 1932 70 1998 260
rect 2044 17 2094 226
rect 2231 364 2281 649
rect 2232 17 2282 226
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 223 390 257 424
rect 991 390 1025 424
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 0 616 50 617
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 979 424 1037 430
rect 979 421 991 424
rect 257 393 991 421
rect 257 390 269 393
rect 211 384 269 390
rect 979 390 991 393
rect 1025 421 1037 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1025 393 1567 421
rect 1025 390 1037 393
rect 979 384 1037 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 49 50 50
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
rlabel locali s 25 200 99 434 6 D
port 1 nsew signal input
rlabel locali s 2130 70 2196 596 6 Q
port 2 nsew signal output
rlabel metal1 s 1555 421 1613 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 384 1613 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 979 421 1037 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 979 384 1037 393 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 421 269 430 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 393 1613 421 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 211 384 269 393 6 RESET_B
port 3 nsew signal input
rlabel locali s 409 346 455 356 6 CLK
port 4 nsew clock input
rlabel locali s 359 264 455 346 6 CLK
port 4 nsew clock input
rlabel metal1 s 0 -49 2304 49 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 617 2304 715 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2943810
string GDS_START 2926420
<< end >>
