magic
tech sky130A
magscale 1 2
timestamp 1604502735
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 17 354 271 649
rect 17 216 127 320
rect 161 250 271 354
rect 17 17 271 216
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 683 288 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 0 617 288 649
rect 0 17 288 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -49 288 -17
<< labels >>
rlabel metal1 s 0 -49 288 49 8 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 617 288 715 6 VPWR
port 2 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 288 666
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 3449026
string GDS_START 3446226
<< end >>
