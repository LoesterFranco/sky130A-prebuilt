magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 103 333 179 493
rect 307 333 373 493
rect 103 299 389 333
rect 22 199 79 265
rect 119 199 215 265
rect 249 199 321 265
rect 119 60 172 199
rect 249 165 283 199
rect 355 165 389 299
rect 435 199 528 333
rect 206 60 283 165
rect 334 51 483 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 299 69 527
rect 223 367 257 527
rect 423 367 479 527
rect 18 17 85 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 435 199 528 333 6 A
port 1 nsew signal input
rlabel locali s 249 199 321 265 6 B
port 2 nsew signal input
rlabel locali s 249 165 283 199 6 B
port 2 nsew signal input
rlabel locali s 206 60 283 165 6 B
port 2 nsew signal input
rlabel locali s 119 199 215 265 6 C
port 3 nsew signal input
rlabel locali s 119 60 172 199 6 C
port 3 nsew signal input
rlabel locali s 22 199 79 265 6 D
port 4 nsew signal input
rlabel locali s 355 165 389 299 6 Y
port 5 nsew signal output
rlabel locali s 334 51 483 165 6 Y
port 5 nsew signal output
rlabel locali s 307 333 373 493 6 Y
port 5 nsew signal output
rlabel locali s 103 333 179 493 6 Y
port 5 nsew signal output
rlabel locali s 103 299 389 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 552 48 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2293008
string GDS_START 2287516
<< end >>
