magic
tech sky130A
magscale 1 2
timestamp 1599588227
<< locali >>
rect 227 401 293 493
rect 457 401 523 493
rect 227 367 523 401
rect 91 199 170 265
rect 291 127 357 367
rect 468 299 523 367
rect 581 255 619 331
rect 422 215 619 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 22 333 82 372
rect 126 367 177 527
rect 345 435 420 527
rect 569 367 603 527
rect 22 299 238 333
rect 22 168 56 299
rect 204 199 238 299
rect 22 102 69 168
rect 119 17 153 155
rect 391 139 619 181
rect 391 93 441 139
rect 207 51 441 93
rect 485 17 519 105
rect 553 51 619 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 91 199 170 265 6 A_N
port 1 nsew signal input
rlabel locali s 581 255 619 331 6 B
port 2 nsew signal input
rlabel locali s 422 215 619 255 6 B
port 2 nsew signal input
rlabel locali s 468 299 523 367 6 Y
port 3 nsew signal output
rlabel locali s 457 401 523 493 6 Y
port 3 nsew signal output
rlabel locali s 291 127 357 367 6 Y
port 3 nsew signal output
rlabel locali s 227 401 293 493 6 Y
port 3 nsew signal output
rlabel locali s 227 367 523 401 6 Y
port 3 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2228600
string GDS_START 2222406
<< end >>
