magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 828 561
rect 18 299 69 527
rect 18 17 69 177
rect 103 59 169 485
rect 232 367 276 527
rect 425 451 491 527
rect 299 199 342 265
rect 203 17 269 93
rect 379 121 433 265
rect 488 199 535 265
rect 579 199 647 265
rect 739 199 801 265
rect 488 121 524 199
rect 644 17 710 97
rect 0 -17 828 17
<< obsli1 >>
rect 318 401 368 493
rect 543 401 605 493
rect 318 367 605 401
rect 759 333 793 493
rect 203 299 793 333
rect 203 165 237 299
rect 203 131 339 165
rect 305 85 339 131
rect 558 131 793 165
rect 558 85 592 131
rect 305 51 592 85
rect 759 51 793 131
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 488 199 535 265 6 A1
port 1 nsew signal input
rlabel locali s 488 121 524 199 6 A1
port 1 nsew signal input
rlabel locali s 379 121 433 265 6 A2
port 2 nsew signal input
rlabel locali s 299 199 342 265 6 A3
port 3 nsew signal input
rlabel locali s 579 199 647 265 6 B1
port 4 nsew signal input
rlabel locali s 739 199 801 265 6 C1
port 5 nsew signal input
rlabel locali s 103 59 169 485 6 X
port 6 nsew signal output
rlabel locali s 644 17 710 97 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 203 17 269 93 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 18 17 69 177 6 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 0 -17 828 17 8 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel locali s 425 451 491 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 232 367 276 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 18 299 69 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 828 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3519014
string GDS_START 3511694
<< end >>
