magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 559 47 589 177
rect 757 47 787 177
rect 841 47 871 177
rect 945 47 975 177
rect 1039 47 1069 177
rect 1123 47 1153 177
rect 1217 47 1247 177
rect 1311 47 1341 177
rect 1415 47 1445 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
<< ndiff >>
rect 27 163 89 177
rect 27 129 35 163
rect 69 129 89 163
rect 27 95 89 129
rect 27 61 35 95
rect 69 61 89 95
rect 27 47 89 61
rect 119 163 173 177
rect 119 129 129 163
rect 163 129 173 163
rect 119 95 173 129
rect 119 61 129 95
rect 163 61 173 95
rect 119 47 173 61
rect 203 163 277 177
rect 203 129 223 163
rect 257 129 277 163
rect 203 47 277 129
rect 307 95 371 177
rect 307 61 317 95
rect 351 61 371 95
rect 307 47 371 61
rect 401 95 455 177
rect 401 61 411 95
rect 445 61 455 95
rect 401 47 455 61
rect 485 163 559 177
rect 485 129 505 163
rect 539 129 559 163
rect 485 95 559 129
rect 485 61 505 95
rect 539 61 559 95
rect 485 47 559 61
rect 589 95 757 177
rect 589 61 599 95
rect 633 61 703 95
rect 737 61 757 95
rect 589 47 757 61
rect 787 163 841 177
rect 787 129 797 163
rect 831 129 841 163
rect 787 95 841 129
rect 787 61 797 95
rect 831 61 841 95
rect 787 47 841 61
rect 871 95 945 177
rect 871 61 891 95
rect 925 61 945 95
rect 871 47 945 61
rect 975 163 1039 177
rect 975 129 985 163
rect 1019 129 1039 163
rect 975 95 1039 129
rect 975 61 985 95
rect 1019 61 1039 95
rect 975 47 1039 61
rect 1069 163 1123 177
rect 1069 129 1079 163
rect 1113 129 1123 163
rect 1069 95 1123 129
rect 1069 61 1079 95
rect 1113 61 1123 95
rect 1069 47 1123 61
rect 1153 163 1217 177
rect 1153 129 1173 163
rect 1207 129 1217 163
rect 1153 95 1217 129
rect 1153 61 1173 95
rect 1207 61 1217 95
rect 1153 47 1217 61
rect 1247 95 1311 177
rect 1247 61 1267 95
rect 1301 61 1311 95
rect 1247 47 1311 61
rect 1341 163 1415 177
rect 1341 129 1361 163
rect 1395 129 1415 163
rect 1341 95 1415 129
rect 1341 61 1361 95
rect 1395 61 1415 95
rect 1341 47 1415 61
rect 1445 95 1497 177
rect 1445 61 1455 95
rect 1489 61 1497 95
rect 1445 47 1497 61
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 297 175 443
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 297 269 375
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 297 363 443
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 341 457 375
rect 399 307 411 341
rect 445 307 457 341
rect 399 297 457 307
rect 493 409 551 497
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 477 641 497
rect 587 443 599 477
rect 633 443 641 477
rect 587 297 641 443
rect 695 485 749 497
rect 695 451 703 485
rect 737 451 749 485
rect 695 297 749 451
rect 785 477 843 497
rect 785 443 797 477
rect 831 443 843 477
rect 785 297 843 443
rect 879 409 937 497
rect 879 375 891 409
rect 925 375 937 409
rect 879 297 937 375
rect 973 477 1031 497
rect 973 443 985 477
rect 1019 443 1031 477
rect 973 409 1031 443
rect 973 375 985 409
rect 1019 375 1031 409
rect 973 297 1031 375
rect 1067 477 1125 497
rect 1067 443 1079 477
rect 1113 443 1125 477
rect 1067 409 1125 443
rect 1067 375 1079 409
rect 1113 375 1125 409
rect 1067 297 1125 375
rect 1161 477 1219 497
rect 1161 443 1173 477
rect 1207 443 1219 477
rect 1161 409 1219 443
rect 1161 375 1173 409
rect 1207 375 1219 409
rect 1161 297 1219 375
rect 1255 483 1313 497
rect 1255 449 1267 483
rect 1301 449 1313 483
rect 1255 297 1313 449
rect 1349 477 1407 497
rect 1349 443 1361 477
rect 1395 443 1407 477
rect 1349 409 1407 443
rect 1349 375 1361 409
rect 1395 375 1407 409
rect 1349 341 1407 375
rect 1349 307 1361 341
rect 1395 307 1407 341
rect 1349 297 1407 307
rect 1443 483 1497 497
rect 1443 449 1455 483
rect 1489 449 1497 483
rect 1443 415 1497 449
rect 1443 381 1455 415
rect 1489 381 1497 415
rect 1443 297 1497 381
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 129 129 163 163
rect 129 61 163 95
rect 223 129 257 163
rect 317 61 351 95
rect 411 61 445 95
rect 505 129 539 163
rect 505 61 539 95
rect 599 61 633 95
rect 703 61 737 95
rect 797 129 831 163
rect 797 61 831 95
rect 891 61 925 95
rect 985 129 1019 163
rect 985 61 1019 95
rect 1079 129 1113 163
rect 1079 61 1113 95
rect 1173 129 1207 163
rect 1173 61 1207 95
rect 1267 61 1301 95
rect 1361 129 1395 163
rect 1361 61 1395 95
rect 1455 61 1489 95
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 443 163 477
rect 223 443 257 477
rect 223 375 257 409
rect 317 443 351 477
rect 411 443 445 477
rect 411 375 445 409
rect 411 307 445 341
rect 505 375 539 409
rect 505 307 539 341
rect 599 443 633 477
rect 703 451 737 485
rect 797 443 831 477
rect 891 375 925 409
rect 985 443 1019 477
rect 985 375 1019 409
rect 1079 443 1113 477
rect 1079 375 1113 409
rect 1173 443 1207 477
rect 1173 375 1207 409
rect 1267 449 1301 483
rect 1361 443 1395 477
rect 1361 375 1395 409
rect 1361 307 1395 341
rect 1455 449 1489 483
rect 1455 381 1489 415
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 79 265 119 282
rect 55 249 119 265
rect 55 215 65 249
rect 99 215 119 249
rect 55 199 119 215
rect 89 177 119 199
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 747 265 787 282
rect 841 265 881 282
rect 935 265 975 282
rect 1029 265 1069 282
rect 1123 265 1163 282
rect 1217 265 1257 282
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 173 249 307 265
rect 173 215 223 249
rect 257 215 307 249
rect 173 199 307 215
rect 349 249 413 265
rect 349 215 359 249
rect 393 215 413 249
rect 349 199 413 215
rect 455 249 649 265
rect 455 215 599 249
rect 633 215 649 249
rect 455 199 649 215
rect 723 249 799 265
rect 723 215 739 249
rect 773 215 799 249
rect 723 199 799 215
rect 841 249 975 265
rect 841 215 857 249
rect 891 215 925 249
rect 959 215 975 249
rect 841 199 975 215
rect 1017 249 1081 265
rect 1017 215 1033 249
rect 1067 215 1081 249
rect 1017 199 1081 215
rect 1123 249 1445 265
rect 1123 215 1199 249
rect 1233 215 1277 249
rect 1311 215 1355 249
rect 1389 215 1445 249
rect 1123 199 1445 215
rect 173 177 203 199
rect 277 177 307 199
rect 371 177 401 199
rect 455 177 485 199
rect 559 177 589 199
rect 757 177 787 199
rect 841 177 871 199
rect 945 177 975 199
rect 1039 177 1069 199
rect 1123 177 1153 199
rect 1217 177 1247 199
rect 1311 177 1341 199
rect 1415 177 1445 199
rect 89 21 119 47
rect 173 21 203 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 559 21 589 47
rect 757 21 787 47
rect 841 21 871 47
rect 945 21 975 47
rect 1039 21 1069 47
rect 1123 21 1153 47
rect 1217 21 1247 47
rect 1311 21 1341 47
rect 1415 21 1445 47
<< polycont >>
rect 65 215 99 249
rect 223 215 257 249
rect 359 215 393 249
rect 599 215 633 249
rect 739 215 773 249
rect 857 215 891 249
rect 925 215 959 249
rect 1033 215 1067 249
rect 1199 215 1233 249
rect 1277 215 1311 249
rect 1355 215 1389 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 27 477 77 493
rect 27 443 35 477
rect 69 443 77 477
rect 27 409 77 443
rect 121 477 171 527
rect 121 443 129 477
rect 163 443 171 477
rect 121 425 171 443
rect 215 477 265 493
rect 215 443 223 477
rect 257 443 265 477
rect 27 375 35 409
rect 69 391 77 409
rect 215 409 265 443
rect 309 477 359 527
rect 309 443 317 477
rect 351 443 359 477
rect 309 425 359 443
rect 403 477 641 493
rect 403 443 411 477
rect 445 459 599 477
rect 445 443 453 459
rect 215 391 223 409
rect 69 375 223 391
rect 257 391 265 409
rect 403 409 453 443
rect 591 443 599 459
rect 633 443 641 477
rect 591 427 641 443
rect 695 485 745 527
rect 695 451 703 485
rect 737 451 745 485
rect 695 427 745 451
rect 789 477 1027 493
rect 789 443 797 477
rect 831 459 985 477
rect 831 443 839 459
rect 789 427 839 443
rect 977 443 985 459
rect 1019 443 1027 477
rect 403 391 411 409
rect 257 375 411 391
rect 445 375 453 409
rect 27 357 453 375
rect 411 341 453 357
rect 17 289 367 323
rect 445 307 453 341
rect 411 291 453 307
rect 497 409 547 425
rect 497 375 505 409
rect 539 393 547 409
rect 883 409 933 425
rect 883 393 891 409
rect 539 375 574 393
rect 497 341 574 375
rect 497 307 505 341
rect 539 323 574 341
rect 687 375 891 393
rect 925 375 933 409
rect 687 357 933 375
rect 977 409 1027 443
rect 977 375 985 409
rect 1019 375 1027 409
rect 977 357 1027 375
rect 1071 477 1121 527
rect 1071 443 1079 477
rect 1113 443 1121 477
rect 1071 409 1121 443
rect 1071 375 1079 409
rect 1113 375 1121 409
rect 1071 359 1121 375
rect 1165 477 1215 493
rect 1165 443 1173 477
rect 1207 443 1215 477
rect 1165 409 1215 443
rect 1259 483 1309 527
rect 1259 449 1267 483
rect 1301 449 1309 483
rect 1259 433 1309 449
rect 1353 477 1403 493
rect 1353 443 1361 477
rect 1395 443 1403 477
rect 1165 375 1173 409
rect 1207 391 1215 409
rect 1353 409 1403 443
rect 1353 391 1361 409
rect 1207 375 1361 391
rect 1395 375 1403 409
rect 1165 357 1403 375
rect 1447 483 1497 527
rect 1447 449 1455 483
rect 1489 449 1497 483
rect 1447 415 1497 449
rect 1447 381 1455 415
rect 1489 381 1497 415
rect 1447 365 1497 381
rect 687 333 721 357
rect 539 307 540 323
rect 17 249 125 289
rect 17 215 65 249
rect 99 215 125 249
rect 171 249 289 255
rect 171 215 223 249
rect 257 215 289 249
rect 333 249 367 289
rect 497 289 540 307
rect 497 283 574 289
rect 651 299 721 333
rect 1353 341 1403 357
rect 333 215 359 249
rect 393 215 419 249
rect 497 181 539 283
rect 651 249 689 299
rect 755 289 1093 323
rect 755 265 801 289
rect 573 215 599 249
rect 633 215 689 249
rect 723 249 801 265
rect 723 215 739 249
rect 773 215 801 249
rect 841 249 983 255
rect 841 215 857 249
rect 891 215 925 249
rect 959 215 983 249
rect 1017 249 1093 289
rect 1017 215 1033 249
rect 1067 215 1093 249
rect 1127 289 1146 323
rect 1180 289 1202 323
rect 1127 249 1202 289
rect 1353 307 1361 341
rect 1395 331 1403 341
rect 1395 307 1535 331
rect 1353 283 1535 307
rect 1127 215 1199 249
rect 1233 215 1277 249
rect 1311 215 1355 249
rect 1389 215 1418 249
rect 651 181 689 215
rect 1462 181 1535 283
rect 35 163 69 179
rect 35 95 69 129
rect 35 17 69 61
rect 103 163 163 181
rect 103 129 129 163
rect 197 163 555 181
rect 197 129 223 163
rect 257 147 505 163
rect 257 129 274 147
rect 479 129 505 147
rect 539 129 555 163
rect 651 163 1035 181
rect 651 145 797 163
rect 103 95 163 129
rect 411 95 445 111
rect 103 61 129 95
rect 163 61 317 95
rect 351 61 367 95
rect 103 51 367 61
rect 411 17 445 61
rect 479 95 555 129
rect 771 129 797 145
rect 831 145 985 163
rect 831 129 847 145
rect 479 61 505 95
rect 539 61 555 95
rect 479 51 555 61
rect 599 95 737 111
rect 633 61 703 95
rect 599 17 737 61
rect 771 95 847 129
rect 959 129 985 145
rect 1019 129 1035 163
rect 771 61 797 95
rect 831 61 847 95
rect 771 51 847 61
rect 891 95 925 111
rect 891 17 925 61
rect 959 95 1035 129
rect 959 61 985 95
rect 1019 61 1035 95
rect 959 51 1035 61
rect 1079 163 1113 179
rect 1079 95 1113 129
rect 1079 17 1113 61
rect 1147 163 1535 181
rect 1147 129 1173 163
rect 1207 145 1361 163
rect 1207 129 1223 145
rect 1147 95 1223 129
rect 1335 129 1361 145
rect 1395 145 1535 163
rect 1395 129 1411 145
rect 1147 61 1173 95
rect 1207 61 1223 95
rect 1147 55 1223 61
rect 1267 95 1301 111
rect 1267 17 1301 61
rect 1335 95 1411 129
rect 1335 61 1361 95
rect 1395 61 1411 95
rect 1335 55 1411 61
rect 1455 95 1489 111
rect 1455 17 1489 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 540 289 574 323
rect 1146 289 1180 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 528 323 596 329
rect 528 289 540 323
rect 574 320 596 323
rect 1134 323 1192 329
rect 1134 320 1146 323
rect 574 292 1146 320
rect 574 289 596 292
rect 528 283 596 289
rect 1134 289 1146 292
rect 1180 289 1192 323
rect 1134 283 1192 289
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel corelocali s 1501 221 1535 255 0 FreeSans 400 180 0 0 X
port 9 nsew
flabel corelocali s 30 221 64 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel corelocali s 212 221 246 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel corelocali s 1501 289 1535 323 0 FreeSans 400 180 0 0 X
port 9 nsew
flabel corelocali s 1041 221 1075 255 0 FreeSans 400 180 0 0 A1_N
port 1 nsew
flabel corelocali s 857 221 891 255 0 FreeSans 400 180 0 0 A2_N
port 2 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1332082
string GDS_START 1320070
<< end >>
