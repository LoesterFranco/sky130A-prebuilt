magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 559 47 589 177
rect 653 47 683 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 561 297 597 497
rect 655 297 691 497
<< ndiff >>
rect 27 119 89 177
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 161 183 177
rect 119 127 129 161
rect 163 127 183 161
rect 119 47 183 127
rect 213 93 277 177
rect 213 59 223 93
rect 257 59 277 93
rect 213 47 277 59
rect 307 161 371 177
rect 307 127 317 161
rect 351 127 371 161
rect 307 47 371 127
rect 401 93 453 177
rect 401 59 411 93
rect 445 59 453 93
rect 401 47 453 59
rect 507 93 559 177
rect 507 59 515 93
rect 549 59 559 93
rect 507 47 559 59
rect 589 161 653 177
rect 589 127 609 161
rect 643 127 653 161
rect 589 47 653 127
rect 683 161 755 177
rect 683 127 709 161
rect 743 127 755 161
rect 683 93 755 127
rect 683 59 709 93
rect 743 59 755 93
rect 683 47 755 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 453 497
rect 399 451 411 485
rect 445 451 453 485
rect 399 417 453 451
rect 399 383 411 417
rect 445 383 453 417
rect 399 297 453 383
rect 507 485 561 497
rect 507 451 515 485
rect 549 451 561 485
rect 507 417 561 451
rect 507 383 515 417
rect 549 383 561 417
rect 507 297 561 383
rect 597 485 655 497
rect 597 451 609 485
rect 643 451 655 485
rect 597 417 655 451
rect 597 383 609 417
rect 643 383 655 417
rect 597 349 655 383
rect 597 315 609 349
rect 643 315 655 349
rect 597 297 655 315
rect 691 485 755 497
rect 691 451 709 485
rect 743 451 755 485
rect 691 417 755 451
rect 691 383 709 417
rect 743 383 755 417
rect 691 349 755 383
rect 691 315 709 349
rect 743 315 755 349
rect 691 297 755 315
<< ndiffc >>
rect 35 85 69 119
rect 129 127 163 161
rect 223 59 257 93
rect 317 127 351 161
rect 411 59 445 93
rect 515 59 549 93
rect 609 127 643 161
rect 709 127 743 161
rect 709 59 743 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 515 451 549 485
rect 515 383 549 417
rect 609 451 643 485
rect 609 383 643 417
rect 609 315 643 349
rect 709 451 743 485
rect 709 383 743 417
rect 709 315 743 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 561 497 597 523
rect 655 497 691 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 561 282 597 297
rect 655 282 691 297
rect 79 265 119 282
rect 173 265 213 282
rect 22 249 213 265
rect 267 261 307 282
rect 361 261 401 282
rect 559 261 599 282
rect 653 263 693 282
rect 653 261 729 263
rect 22 215 32 249
rect 66 215 213 249
rect 22 199 213 215
rect 255 249 437 261
rect 255 215 271 249
rect 305 215 377 249
rect 411 215 437 249
rect 255 203 437 215
rect 559 249 729 261
rect 559 215 575 249
rect 609 215 669 249
rect 703 215 729 249
rect 559 203 729 215
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 203
rect 371 177 401 203
rect 559 177 589 203
rect 653 202 729 203
rect 653 177 683 202
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 559 21 589 47
rect 653 21 683 47
<< polycont >>
rect 32 215 66 249
rect 271 215 305 249
rect 377 215 411 249
rect 575 215 609 249
rect 669 215 703 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 549 527
rect 445 451 515 485
rect 411 417 549 451
rect 445 383 515 417
rect 411 367 549 383
rect 583 485 659 493
rect 583 451 609 485
rect 643 451 659 485
rect 583 417 659 451
rect 583 383 609 417
rect 643 383 659 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 583 349 659 383
rect 583 333 609 349
rect 351 315 609 333
rect 643 315 659 349
rect 103 289 659 315
rect 703 485 779 527
rect 703 451 709 485
rect 743 451 779 485
rect 703 417 779 451
rect 703 383 709 417
rect 743 383 779 417
rect 703 349 779 383
rect 703 315 709 349
rect 743 315 779 349
rect 703 289 779 315
rect 18 249 66 265
rect 18 215 32 249
rect 18 199 66 215
rect 103 161 179 289
rect 234 249 523 255
rect 234 215 271 249
rect 305 215 377 249
rect 411 215 523 249
rect 557 249 800 255
rect 557 215 575 249
rect 609 215 669 249
rect 703 215 800 249
rect 18 119 69 157
rect 103 127 129 161
rect 163 127 179 161
rect 291 161 659 181
rect 291 127 317 161
rect 351 127 609 161
rect 643 127 659 161
rect 703 161 779 177
rect 703 127 709 161
rect 743 127 779 161
rect 18 85 35 119
rect 703 93 779 127
rect 69 85 223 93
rect 18 59 223 85
rect 257 59 411 93
rect 445 59 461 93
rect 499 59 515 93
rect 549 59 565 93
rect 499 17 565 59
rect 703 59 709 93
rect 743 59 779 93
rect 703 17 779 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel corelocali s 30 221 64 255 0 FreeSans 250 0 0 0 A
port 1 nsew
flabel corelocali s 132 153 166 187 0 FreeSans 250 0 0 0 Y
port 8 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 250 0 0 0 Y
port 8 nsew
flabel corelocali s 132 289 166 323 0 FreeSans 250 0 0 0 Y
port 8 nsew
flabel corelocali s 480 221 514 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 302 221 336 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 396 221 430 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel corelocali s 676 221 710 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 585 221 619 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel corelocali s 764 221 798 255 0 FreeSans 250 0 0 0 C
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
rlabel comment s 0 0 0 0 4 nand3_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2250328
string GDS_START 2242750
<< end >>
