magic
tech sky130A
magscale 1 2
timestamp 1604502701
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 0 0 1440 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 286 368 316 592
rect 376 368 406 592
rect 588 392 618 592
rect 692 392 722 592
rect 812 392 842 592
rect 922 392 952 592
rect 1012 392 1042 592
rect 1124 392 1154 592
rect 1224 392 1254 592
rect 1324 392 1354 592
<< nmoslvt >>
rect 89 74 119 222
rect 184 74 214 222
rect 270 74 300 222
rect 361 74 391 222
rect 559 74 589 202
rect 659 74 689 202
rect 745 74 775 202
rect 845 74 875 202
rect 1057 74 1087 202
rect 1143 74 1173 202
rect 1229 74 1259 202
rect 1315 74 1345 202
<< ndiff >>
rect 27 210 89 222
rect 27 176 39 210
rect 73 176 89 210
rect 27 120 89 176
rect 27 86 39 120
rect 73 86 89 120
rect 27 74 89 86
rect 119 210 184 222
rect 119 176 139 210
rect 173 176 184 210
rect 119 120 184 176
rect 119 86 139 120
rect 173 86 184 120
rect 119 74 184 86
rect 214 130 270 222
rect 214 96 225 130
rect 259 96 270 130
rect 214 74 270 96
rect 300 184 361 222
rect 300 150 311 184
rect 345 150 361 184
rect 300 116 361 150
rect 300 82 311 116
rect 345 82 361 116
rect 300 74 361 82
rect 391 188 448 222
rect 391 154 402 188
rect 436 154 448 188
rect 391 120 448 154
rect 391 86 402 120
rect 436 86 448 120
rect 391 74 448 86
rect 502 190 559 202
rect 502 156 514 190
rect 548 156 559 190
rect 502 120 559 156
rect 502 86 514 120
rect 548 86 559 120
rect 502 74 559 86
rect 589 184 659 202
rect 589 150 600 184
rect 634 150 659 184
rect 589 116 659 150
rect 589 82 600 116
rect 634 82 659 116
rect 589 74 659 82
rect 689 190 745 202
rect 689 156 700 190
rect 734 156 745 190
rect 689 120 745 156
rect 689 86 700 120
rect 734 86 745 120
rect 689 74 745 86
rect 775 184 845 202
rect 775 150 800 184
rect 834 150 845 184
rect 775 116 845 150
rect 775 82 800 116
rect 834 82 845 116
rect 775 74 845 82
rect 875 169 946 202
rect 875 135 900 169
rect 934 135 946 169
rect 875 74 946 135
rect 1000 169 1057 202
rect 1000 135 1012 169
rect 1046 135 1057 169
rect 1000 74 1057 135
rect 1087 184 1143 202
rect 1087 150 1098 184
rect 1132 150 1143 184
rect 1087 116 1143 150
rect 1087 82 1098 116
rect 1132 82 1143 116
rect 1087 74 1143 82
rect 1173 190 1229 202
rect 1173 156 1184 190
rect 1218 156 1229 190
rect 1173 120 1229 156
rect 1173 86 1184 120
rect 1218 86 1229 120
rect 1173 74 1229 86
rect 1259 184 1315 202
rect 1259 150 1270 184
rect 1304 150 1315 184
rect 1259 116 1315 150
rect 1259 82 1270 116
rect 1304 82 1315 116
rect 1259 74 1315 82
rect 1345 190 1402 202
rect 1345 156 1356 190
rect 1390 156 1402 190
rect 1345 120 1402 156
rect 1345 86 1356 120
rect 1390 86 1402 120
rect 1345 74 1402 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 497 176 546
rect 116 463 129 497
rect 163 463 176 497
rect 116 414 176 463
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 582 286 592
rect 206 548 229 582
rect 263 548 286 582
rect 206 514 286 548
rect 206 480 229 514
rect 263 480 286 514
rect 206 446 286 480
rect 206 412 229 446
rect 263 412 286 446
rect 206 368 286 412
rect 316 580 376 592
rect 316 546 329 580
rect 363 546 376 580
rect 316 497 376 546
rect 316 463 329 497
rect 363 463 376 497
rect 316 414 376 463
rect 316 380 329 414
rect 363 380 376 414
rect 316 368 376 380
rect 406 580 475 592
rect 406 546 429 580
rect 463 546 475 580
rect 406 497 475 546
rect 406 463 429 497
rect 463 463 475 497
rect 406 414 475 463
rect 406 380 429 414
rect 463 380 475 414
rect 529 580 588 592
rect 529 546 541 580
rect 575 546 588 580
rect 529 512 588 546
rect 529 478 541 512
rect 575 478 588 512
rect 529 444 588 478
rect 529 410 541 444
rect 575 410 588 444
rect 529 392 588 410
rect 618 519 692 592
rect 618 485 643 519
rect 677 485 692 519
rect 618 434 692 485
rect 618 400 643 434
rect 677 400 692 434
rect 618 392 692 400
rect 722 580 812 592
rect 722 546 765 580
rect 799 546 812 580
rect 722 510 812 546
rect 722 476 765 510
rect 799 476 812 510
rect 722 440 812 476
rect 722 406 765 440
rect 799 406 812 440
rect 722 392 812 406
rect 842 580 922 592
rect 842 546 865 580
rect 899 546 922 580
rect 842 502 922 546
rect 842 468 865 502
rect 899 468 922 502
rect 842 392 922 468
rect 952 580 1012 592
rect 952 546 965 580
rect 999 546 1012 580
rect 952 510 1012 546
rect 952 476 965 510
rect 999 476 1012 510
rect 952 440 1012 476
rect 952 406 965 440
rect 999 406 1012 440
rect 952 392 1012 406
rect 1042 580 1124 592
rect 1042 546 1065 580
rect 1099 546 1124 580
rect 1042 502 1124 546
rect 1042 468 1065 502
rect 1099 468 1124 502
rect 1042 392 1124 468
rect 1154 580 1224 592
rect 1154 546 1167 580
rect 1201 546 1224 580
rect 1154 510 1224 546
rect 1154 476 1167 510
rect 1201 476 1224 510
rect 1154 440 1224 476
rect 1154 406 1167 440
rect 1201 406 1224 440
rect 1154 392 1224 406
rect 1254 580 1324 592
rect 1254 546 1267 580
rect 1301 546 1324 580
rect 1254 502 1324 546
rect 1254 468 1267 502
rect 1301 468 1324 502
rect 1254 392 1324 468
rect 1354 580 1413 592
rect 1354 546 1367 580
rect 1401 546 1413 580
rect 1354 510 1413 546
rect 1354 476 1367 510
rect 1401 476 1413 510
rect 1354 440 1413 476
rect 1354 406 1367 440
rect 1401 406 1413 440
rect 1354 392 1413 406
rect 406 368 475 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 225 96 259 130
rect 311 150 345 184
rect 311 82 345 116
rect 402 154 436 188
rect 402 86 436 120
rect 514 156 548 190
rect 514 86 548 120
rect 600 150 634 184
rect 600 82 634 116
rect 700 156 734 190
rect 700 86 734 120
rect 800 150 834 184
rect 800 82 834 116
rect 900 135 934 169
rect 1012 135 1046 169
rect 1098 150 1132 184
rect 1098 82 1132 116
rect 1184 156 1218 190
rect 1184 86 1218 120
rect 1270 150 1304 184
rect 1270 82 1304 116
rect 1356 156 1390 190
rect 1356 86 1390 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 229 548 263 582
rect 229 480 263 514
rect 229 412 263 446
rect 329 546 363 580
rect 329 463 363 497
rect 329 380 363 414
rect 429 546 463 580
rect 429 463 463 497
rect 429 380 463 414
rect 541 546 575 580
rect 541 478 575 512
rect 541 410 575 444
rect 643 485 677 519
rect 643 400 677 434
rect 765 546 799 580
rect 765 476 799 510
rect 765 406 799 440
rect 865 546 899 580
rect 865 468 899 502
rect 965 546 999 580
rect 965 476 999 510
rect 965 406 999 440
rect 1065 546 1099 580
rect 1065 468 1099 502
rect 1167 546 1201 580
rect 1167 476 1201 510
rect 1167 406 1201 440
rect 1267 546 1301 580
rect 1267 468 1301 502
rect 1367 546 1401 580
rect 1367 476 1401 510
rect 1367 406 1401 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 286 592 316 618
rect 376 592 406 618
rect 588 592 618 618
rect 692 592 722 618
rect 812 592 842 618
rect 922 592 952 618
rect 1012 592 1042 618
rect 1124 592 1154 618
rect 1224 592 1254 618
rect 1324 592 1354 618
rect 588 377 618 392
rect 692 377 722 392
rect 812 377 842 392
rect 922 377 952 392
rect 1012 377 1042 392
rect 1124 377 1154 392
rect 1224 377 1254 392
rect 1324 377 1354 392
rect 86 353 116 368
rect 176 353 206 368
rect 286 353 316 368
rect 376 353 406 368
rect 585 360 621 377
rect 689 360 725 377
rect 83 310 119 353
rect 173 310 209 353
rect 283 310 319 353
rect 373 310 409 353
rect 513 344 725 360
rect 513 310 529 344
rect 563 310 597 344
rect 631 330 725 344
rect 809 356 845 377
rect 919 356 955 377
rect 809 340 955 356
rect 631 310 689 330
rect 83 294 467 310
rect 513 294 689 310
rect 83 274 213 294
rect 89 260 213 274
rect 247 260 281 294
rect 315 260 349 294
rect 383 260 417 294
rect 451 260 467 294
rect 89 244 467 260
rect 89 222 119 244
rect 184 222 214 244
rect 270 222 300 244
rect 361 222 391 244
rect 559 202 589 294
rect 659 202 689 294
rect 809 306 825 340
rect 859 306 893 340
rect 927 306 955 340
rect 1009 356 1045 377
rect 1121 356 1157 377
rect 1221 356 1257 377
rect 1321 356 1357 377
rect 1009 340 1173 356
rect 1009 320 1055 340
rect 809 290 955 306
rect 1015 306 1055 320
rect 1089 306 1123 340
rect 1157 306 1173 340
rect 1015 290 1173 306
rect 1221 340 1357 356
rect 1221 306 1239 340
rect 1273 306 1307 340
rect 1341 306 1357 340
rect 1221 290 1357 306
rect 809 247 875 290
rect 745 217 875 247
rect 1015 247 1045 290
rect 1015 217 1087 247
rect 745 202 775 217
rect 845 202 875 217
rect 1057 202 1087 217
rect 1143 202 1173 290
rect 1229 202 1259 290
rect 1315 202 1345 290
rect 89 48 119 74
rect 184 48 214 74
rect 270 48 300 74
rect 361 48 391 74
rect 559 48 589 74
rect 659 48 689 74
rect 745 48 775 74
rect 845 48 875 74
rect 1057 48 1087 74
rect 1143 48 1173 74
rect 1229 48 1259 74
rect 1315 48 1345 74
<< polycont >>
rect 529 310 563 344
rect 597 310 631 344
rect 213 260 247 294
rect 281 260 315 294
rect 349 260 383 294
rect 417 260 451 294
rect 825 306 859 340
rect 893 306 927 340
rect 1055 306 1089 340
rect 1123 306 1157 340
rect 1239 306 1273 340
rect 1307 306 1341 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 497 179 546
rect 113 463 129 497
rect 163 463 179 497
rect 113 414 179 463
rect 113 380 129 414
rect 163 380 179 414
rect 213 582 279 649
rect 213 548 229 582
rect 263 548 279 582
rect 213 514 279 548
rect 213 480 229 514
rect 263 480 279 514
rect 213 446 279 480
rect 213 412 229 446
rect 263 412 279 446
rect 313 580 379 596
rect 313 546 329 580
rect 363 546 379 580
rect 313 497 379 546
rect 313 463 329 497
rect 363 463 379 497
rect 313 414 379 463
rect 113 378 179 380
rect 313 380 329 414
rect 363 380 379 414
rect 313 378 379 380
rect 113 344 379 378
rect 413 580 479 649
rect 413 546 429 580
rect 463 546 479 580
rect 413 497 479 546
rect 413 463 429 497
rect 463 463 479 497
rect 413 414 479 463
rect 413 380 429 414
rect 463 380 479 414
rect 525 580 815 596
rect 525 546 541 580
rect 575 562 765 580
rect 575 546 591 562
rect 525 512 591 546
rect 749 546 765 562
rect 799 546 815 580
rect 525 478 541 512
rect 575 478 591 512
rect 525 444 591 478
rect 525 410 541 444
rect 575 410 591 444
rect 525 394 591 410
rect 625 519 715 528
rect 625 485 643 519
rect 677 485 715 519
rect 625 434 715 485
rect 625 400 643 434
rect 677 400 715 434
rect 625 394 715 400
rect 413 364 479 380
rect 513 344 647 360
rect 113 310 179 344
rect 513 310 529 344
rect 563 310 597 344
rect 631 310 647 344
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 173 310
rect 213 294 467 310
rect 513 294 647 310
rect 247 260 281 294
rect 315 260 349 294
rect 383 260 417 294
rect 451 260 467 294
rect 681 260 715 394
rect 749 510 815 546
rect 749 476 765 510
rect 799 476 815 510
rect 749 440 815 476
rect 849 580 915 649
rect 849 546 865 580
rect 899 546 915 580
rect 849 502 915 546
rect 849 468 865 502
rect 899 468 915 502
rect 849 458 915 468
rect 949 580 1015 596
rect 949 546 965 580
rect 999 546 1015 580
rect 949 510 1015 546
rect 949 476 965 510
rect 999 476 1015 510
rect 749 406 765 440
rect 799 424 815 440
rect 949 440 1015 476
rect 1049 580 1115 649
rect 1049 546 1065 580
rect 1099 546 1115 580
rect 1049 502 1115 546
rect 1049 468 1065 502
rect 1099 468 1115 502
rect 1049 458 1115 468
rect 1151 580 1217 596
rect 1151 546 1167 580
rect 1201 546 1217 580
rect 1151 510 1217 546
rect 1151 476 1167 510
rect 1201 476 1217 510
rect 949 424 965 440
rect 799 406 965 424
rect 999 424 1015 440
rect 1151 440 1217 476
rect 1251 580 1317 649
rect 1251 546 1267 580
rect 1301 546 1317 580
rect 1251 502 1317 546
rect 1251 468 1267 502
rect 1301 468 1317 502
rect 1251 458 1317 468
rect 1351 580 1417 596
rect 1351 546 1367 580
rect 1401 546 1417 580
rect 1351 510 1417 546
rect 1351 476 1367 510
rect 1401 476 1417 510
rect 1151 424 1167 440
rect 999 406 1167 424
rect 1201 424 1217 440
rect 1351 440 1417 476
rect 1351 424 1367 440
rect 1201 406 1367 424
rect 1401 406 1417 440
rect 749 390 1417 406
rect 793 340 935 356
rect 793 306 825 340
rect 859 306 893 340
rect 927 306 935 340
rect 793 290 935 306
rect 985 340 1173 356
rect 985 306 1055 340
rect 1089 306 1123 340
rect 1157 306 1173 340
rect 985 290 1173 306
rect 1223 340 1415 356
rect 1223 306 1239 340
rect 1273 306 1307 340
rect 1341 306 1415 340
rect 1223 290 1415 306
rect 213 256 718 260
rect 213 244 950 256
rect 379 226 950 244
rect 123 176 139 210
rect 173 184 345 200
rect 173 176 311 184
rect 123 166 311 176
rect 123 120 173 166
rect 123 86 139 120
rect 123 70 173 86
rect 209 130 275 132
rect 209 96 225 130
rect 259 96 275 130
rect 209 17 275 96
rect 311 116 345 150
rect 311 66 345 82
rect 386 188 452 192
rect 386 154 402 188
rect 436 154 452 188
rect 386 120 452 154
rect 386 86 402 120
rect 436 86 452 120
rect 386 17 452 86
rect 498 190 548 226
rect 684 222 950 226
rect 498 156 514 190
rect 498 120 548 156
rect 498 86 514 120
rect 498 70 548 86
rect 584 184 650 192
rect 584 150 600 184
rect 634 150 650 184
rect 584 116 650 150
rect 584 82 600 116
rect 634 82 650 116
rect 584 17 650 82
rect 684 190 750 222
rect 684 156 700 190
rect 734 156 750 190
rect 684 120 750 156
rect 684 86 700 120
rect 734 86 750 120
rect 684 70 750 86
rect 784 184 850 188
rect 784 150 800 184
rect 834 150 850 184
rect 784 116 850 150
rect 884 169 950 222
rect 884 135 900 169
rect 934 135 950 169
rect 884 119 950 135
rect 996 222 1406 256
rect 996 169 1046 222
rect 1184 190 1218 222
rect 996 135 1012 169
rect 996 119 1046 135
rect 1082 184 1148 188
rect 1082 150 1098 184
rect 1132 150 1148 184
rect 784 82 800 116
rect 834 85 850 116
rect 1082 116 1148 150
rect 1082 85 1098 116
rect 834 82 1098 85
rect 1132 82 1148 116
rect 784 51 1148 82
rect 1356 190 1406 222
rect 1184 120 1218 156
rect 1184 70 1218 86
rect 1254 184 1320 188
rect 1254 150 1270 184
rect 1304 150 1320 184
rect 1254 116 1320 150
rect 1254 82 1270 116
rect 1304 82 1320 116
rect 1254 17 1320 82
rect 1390 156 1406 190
rect 1356 120 1406 156
rect 1390 86 1406 120
rect 1356 70 1406 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a31o_4
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nbase s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew
flabel corelocali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew
flabel corelocali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew
flabel corelocali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A3
port 3 nsew
flabel corelocali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew
flabel corelocali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 9 nsew
flabel corelocali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 1440 666
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3802782
string GDS_START 3789944
<< end >>
