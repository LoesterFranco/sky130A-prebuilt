magic
tech sky130A
magscale 1 2
timestamp 1601050047
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 94 424 124 592
rect 338 391 368 591
rect 422 391 452 591
rect 506 391 536 591
rect 623 368 653 592
<< nmoslvt >>
rect 97 74 127 184
rect 296 74 326 184
rect 410 74 440 184
rect 503 74 533 184
rect 654 74 684 222
<< ndiff >>
rect 604 184 654 222
rect 27 146 97 184
rect 27 112 39 146
rect 73 112 97 146
rect 27 74 97 112
rect 127 146 185 184
rect 127 112 139 146
rect 173 112 185 146
rect 127 74 185 112
rect 239 146 296 184
rect 239 112 251 146
rect 285 112 296 146
rect 239 74 296 112
rect 326 120 410 184
rect 326 86 351 120
rect 385 86 410 120
rect 326 74 410 86
rect 440 146 503 184
rect 440 112 451 146
rect 485 112 503 146
rect 440 74 503 112
rect 533 120 654 184
rect 533 86 573 120
rect 607 86 654 120
rect 533 74 654 86
rect 684 210 741 222
rect 684 176 695 210
rect 729 176 741 210
rect 684 120 741 176
rect 684 86 695 120
rect 729 86 741 120
rect 684 74 741 86
<< pdiff >>
rect 27 580 94 592
rect 27 546 39 580
rect 73 546 94 580
rect 27 470 94 546
rect 27 436 39 470
rect 73 436 94 470
rect 27 424 94 436
rect 124 580 185 592
rect 554 591 623 592
rect 124 546 139 580
rect 173 546 185 580
rect 124 470 185 546
rect 124 436 139 470
rect 173 436 185 470
rect 124 424 185 436
rect 279 579 338 591
rect 279 545 291 579
rect 325 545 338 579
rect 279 508 338 545
rect 279 474 291 508
rect 325 474 338 508
rect 279 437 338 474
rect 279 403 291 437
rect 325 403 338 437
rect 279 391 338 403
rect 368 391 422 591
rect 452 391 506 591
rect 536 580 623 591
rect 536 546 566 580
rect 600 546 623 580
rect 536 510 623 546
rect 536 476 566 510
rect 600 476 623 510
rect 536 440 623 476
rect 536 406 566 440
rect 600 406 623 440
rect 536 391 623 406
rect 554 368 623 391
rect 653 580 712 592
rect 653 546 666 580
rect 700 546 712 580
rect 653 497 712 546
rect 653 463 666 497
rect 700 463 712 497
rect 653 414 712 463
rect 653 380 666 414
rect 700 380 712 414
rect 653 368 712 380
<< ndiffc >>
rect 39 112 73 146
rect 139 112 173 146
rect 251 112 285 146
rect 351 86 385 120
rect 451 112 485 146
rect 573 86 607 120
rect 695 176 729 210
rect 695 86 729 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 139 546 173 580
rect 139 436 173 470
rect 291 545 325 579
rect 291 474 325 508
rect 291 403 325 437
rect 566 546 600 580
rect 566 476 600 510
rect 566 406 600 440
rect 666 546 700 580
rect 666 463 700 497
rect 666 380 700 414
<< poly >>
rect 94 592 124 618
rect 338 591 368 617
rect 422 591 452 617
rect 506 591 536 617
rect 623 592 653 618
rect 94 409 124 424
rect 91 356 127 409
rect 338 376 368 391
rect 422 376 452 391
rect 506 376 536 391
rect 55 340 127 356
rect 55 306 71 340
rect 105 306 127 340
rect 55 272 127 306
rect 55 238 71 272
rect 105 238 127 272
rect 175 360 371 376
rect 175 326 191 360
rect 225 346 371 360
rect 225 326 241 346
rect 175 292 241 326
rect 419 304 455 376
rect 503 326 539 376
rect 623 353 653 368
rect 620 326 656 353
rect 503 310 569 326
rect 175 258 191 292
rect 225 272 241 292
rect 383 288 449 304
rect 225 258 326 272
rect 175 242 326 258
rect 55 222 127 238
rect 97 184 127 222
rect 296 184 326 242
rect 383 254 399 288
rect 433 254 449 288
rect 383 238 449 254
rect 503 276 519 310
rect 553 276 569 310
rect 503 260 569 276
rect 617 310 684 326
rect 617 276 633 310
rect 667 276 684 310
rect 617 260 684 276
rect 410 184 440 238
rect 503 184 533 260
rect 654 222 684 260
rect 97 48 127 74
rect 296 48 326 74
rect 410 48 440 74
rect 503 48 533 74
rect 654 48 684 74
<< polycont >>
rect 71 306 105 340
rect 71 238 105 272
rect 191 326 225 360
rect 191 258 225 292
rect 399 254 433 288
rect 519 276 553 310
rect 633 276 667 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 470 89 546
rect 23 436 39 470
rect 73 436 89 470
rect 23 420 89 436
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 470 189 546
rect 123 436 139 470
rect 173 436 189 470
rect 123 420 189 436
rect 155 376 189 420
rect 275 579 341 595
rect 275 545 291 579
rect 325 545 341 579
rect 550 580 616 649
rect 275 508 341 545
rect 275 474 291 508
rect 325 474 341 508
rect 275 437 341 474
rect 275 403 291 437
rect 325 403 341 437
rect 155 360 241 376
rect 25 340 121 356
rect 25 306 71 340
rect 105 306 121 340
rect 25 272 121 306
rect 25 238 71 272
rect 105 238 121 272
rect 25 222 121 238
rect 155 326 191 360
rect 225 326 241 360
rect 155 292 241 326
rect 155 258 191 292
rect 225 258 241 292
rect 155 242 241 258
rect 155 188 189 242
rect 275 204 341 403
rect 383 288 455 578
rect 550 546 566 580
rect 600 546 616 580
rect 550 510 616 546
rect 550 476 566 510
rect 600 476 616 510
rect 550 440 616 476
rect 550 406 566 440
rect 600 406 616 440
rect 550 390 616 406
rect 650 580 751 596
rect 650 546 666 580
rect 700 546 751 580
rect 650 497 751 546
rect 650 463 666 497
rect 700 463 751 497
rect 650 414 751 463
rect 650 380 666 414
rect 700 380 751 414
rect 650 364 751 380
rect 383 254 399 288
rect 433 254 455 288
rect 503 310 569 356
rect 503 276 519 310
rect 553 276 569 310
rect 503 260 569 276
rect 611 310 683 326
rect 611 276 633 310
rect 667 276 683 310
rect 611 260 683 276
rect 383 238 455 254
rect 611 204 645 260
rect 717 226 751 364
rect 23 146 89 188
rect 23 112 39 146
rect 73 112 89 146
rect 23 17 89 112
rect 123 146 189 188
rect 123 112 139 146
rect 173 112 189 146
rect 123 70 189 112
rect 235 170 645 204
rect 679 210 751 226
rect 679 176 695 210
rect 729 176 751 210
rect 235 146 301 170
rect 235 112 251 146
rect 285 112 301 146
rect 435 146 501 170
rect 235 70 301 112
rect 335 120 401 136
rect 335 86 351 120
rect 385 86 401 120
rect 335 17 401 86
rect 435 112 451 146
rect 485 112 501 146
rect 435 70 501 112
rect 535 120 645 136
rect 535 86 573 120
rect 607 86 645 120
rect 535 17 645 86
rect 679 120 751 176
rect 679 86 695 120
rect 729 86 751 120
rect 679 70 751 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or3b_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel corelocali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 390 449 424 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 464 449 498 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 415 538 449 572 0 FreeSans 340 0 0 0 B
port 2 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew
flabel corelocali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 8 nsew
flabel corelocali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 768 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 820256
string GDS_START 813042
<< end >>
