magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 384 370 463 596
rect 215 236 281 336
rect 429 236 463 370
rect 21 51 167 134
rect 368 94 463 236
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 70 438 137 649
rect 171 404 237 600
rect 278 438 344 649
rect 52 370 350 404
rect 52 168 118 370
rect 316 336 350 370
rect 316 270 395 336
rect 268 17 334 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
rlabel locali s 21 51 167 134 6 A
port 1 nsew signal input
rlabel locali s 215 236 281 336 6 B
port 2 nsew signal input
rlabel locali s 429 236 463 370 6 X
port 3 nsew signal output
rlabel locali s 384 370 463 596 6 X
port 3 nsew signal output
rlabel locali s 368 94 463 236 6 X
port 3 nsew signal output
rlabel metal1 s 0 -49 480 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 480 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 3191460
string GDS_START 3186388
<< end >>
