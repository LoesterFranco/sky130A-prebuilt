magic
tech sky130A
magscale 1 2
timestamp 1601050070
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 35 367 69 527
rect 223 367 257 527
rect 411 367 445 527
rect 505 323 539 493
rect 573 367 649 527
rect 693 323 727 493
rect 761 367 837 527
rect 881 323 915 493
rect 949 367 1025 527
rect 1069 323 1103 493
rect 1137 367 1213 527
rect 1257 323 1291 493
rect 1325 367 1401 527
rect 1445 323 1479 493
rect 505 289 1479 323
rect 1513 297 1589 527
rect 27 215 362 255
rect 1042 181 1479 289
rect 505 147 1479 181
rect 19 17 85 113
rect 197 17 273 113
rect 385 17 461 113
rect 505 51 539 147
rect 573 17 649 113
rect 693 51 727 147
rect 761 17 837 113
rect 881 51 915 147
rect 949 17 1025 113
rect 1069 51 1103 147
rect 1137 17 1213 113
rect 1257 51 1291 147
rect 1325 17 1401 113
rect 1445 51 1479 147
rect 1513 17 1589 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< obsli1 >>
rect 103 323 179 493
rect 291 323 367 493
rect 103 289 443 323
rect 408 249 443 289
rect 408 215 993 249
rect 408 181 443 215
rect 129 147 443 181
rect 129 51 163 147
rect 317 52 351 147
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
rlabel locali s 27 215 362 255 6 A
port 1 nsew signal input
rlabel locali s 1445 323 1479 493 6 X
port 2 nsew signal output
rlabel locali s 1445 51 1479 147 6 X
port 2 nsew signal output
rlabel locali s 1257 323 1291 493 6 X
port 2 nsew signal output
rlabel locali s 1257 51 1291 147 6 X
port 2 nsew signal output
rlabel locali s 1069 323 1103 493 6 X
port 2 nsew signal output
rlabel locali s 1069 51 1103 147 6 X
port 2 nsew signal output
rlabel locali s 1042 181 1479 289 6 X
port 2 nsew signal output
rlabel locali s 881 323 915 493 6 X
port 2 nsew signal output
rlabel locali s 881 51 915 147 6 X
port 2 nsew signal output
rlabel locali s 693 323 727 493 6 X
port 2 nsew signal output
rlabel locali s 693 51 727 147 6 X
port 2 nsew signal output
rlabel locali s 505 323 539 493 6 X
port 2 nsew signal output
rlabel locali s 505 289 1479 323 6 X
port 2 nsew signal output
rlabel locali s 505 147 1479 181 6 X
port 2 nsew signal output
rlabel locali s 505 51 539 147 6 X
port 2 nsew signal output
rlabel viali s 1593 -17 1627 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 1501 -17 1535 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 1409 -17 1443 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 1317 -17 1351 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 1225 -17 1259 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 1133 -17 1167 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 1041 -17 1075 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 949 -17 983 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 857 -17 891 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 765 -17 799 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 673 -17 707 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 581 -17 615 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 489 -17 523 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 397 -17 431 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 305 -17 339 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 213 -17 247 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 121 -17 155 17 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 29 -17 63 17 8 VGND
port 3 nsew ground bidirectional
rlabel locali s 1513 17 1589 177 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 1325 17 1401 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 1137 17 1213 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 949 17 1025 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 761 17 837 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 573 17 649 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 385 17 461 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 197 17 273 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 19 17 85 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 0 -17 1656 17 8 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -48 1656 48 8 VGND
port 3 nsew ground bidirectional
rlabel viali s 1593 527 1627 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 1501 527 1535 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 1409 527 1443 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 1317 527 1351 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 1225 527 1259 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 1133 527 1167 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 1041 527 1075 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 949 527 983 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 857 527 891 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 765 527 799 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 673 527 707 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 581 527 615 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 489 527 523 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 397 527 431 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 305 527 339 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 213 527 247 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 121 527 155 561 6 VPWR
port 4 nsew power bidirectional
rlabel viali s 29 527 63 561 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 1513 297 1589 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 1325 367 1401 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 1137 367 1213 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 949 367 1025 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 761 367 837 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 573 367 649 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 411 367 445 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 223 367 257 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 35 367 69 527 6 VPWR
port 4 nsew power bidirectional
rlabel locali s 0 527 1656 561 6 VPWR
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1639512
string GDS_START 1627650
<< end >>
