magic
tech sky130A
magscale 1 2
timestamp 1601050052
<< nwell >>
rect -38 335 2246 704
rect -38 332 645 335
rect 1384 332 2246 335
rect 187 311 645 332
<< pwell >>
rect 0 0 2208 49
<< scnmos >>
rect 90 74 120 158
rect 168 74 198 158
rect 270 74 300 222
rect 480 79 510 227
rect 684 127 714 211
rect 820 127 850 211
rect 892 127 922 211
rect 964 127 994 211
rect 1148 119 1178 267
rect 1236 119 1266 267
rect 1520 119 1550 203
rect 1598 119 1628 203
rect 1706 119 1736 203
rect 1784 119 1814 203
rect 1991 94 2021 204
rect 2093 94 2123 242
<< pmoshvt >>
rect 85 508 115 592
rect 175 508 205 592
rect 276 347 306 547
rect 477 347 507 547
rect 697 463 727 547
rect 787 463 817 547
rect 865 463 895 547
rect 964 463 994 547
rect 1161 392 1191 592
rect 1347 392 1377 592
rect 1517 508 1547 592
rect 1601 508 1631 592
rect 1709 508 1739 592
rect 1799 508 1829 592
rect 1993 424 2023 592
rect 2094 368 2124 592
<< ndiff >>
rect 213 158 270 222
rect 33 131 90 158
rect 33 97 45 131
rect 79 97 90 131
rect 33 74 90 97
rect 120 74 168 158
rect 198 133 270 158
rect 198 99 225 133
rect 259 99 270 133
rect 198 74 270 99
rect 300 202 355 222
rect 300 168 311 202
rect 345 168 355 202
rect 300 120 355 168
rect 300 86 311 120
rect 345 86 355 120
rect 300 74 355 86
rect 409 79 480 227
rect 510 215 577 227
rect 510 181 535 215
rect 569 181 577 215
rect 1098 211 1148 267
rect 510 79 577 181
rect 631 188 684 211
rect 631 154 639 188
rect 673 154 684 188
rect 631 127 684 154
rect 714 188 820 211
rect 714 154 775 188
rect 809 154 820 188
rect 714 127 820 154
rect 850 127 892 211
rect 922 127 964 211
rect 994 127 1148 211
rect 409 77 465 79
rect 409 43 417 77
rect 451 43 465 77
rect 409 31 465 43
rect 1009 124 1148 127
rect 1009 90 1021 124
rect 1055 119 1148 124
rect 1178 244 1236 267
rect 1178 210 1189 244
rect 1223 210 1236 244
rect 1178 169 1236 210
rect 1178 135 1189 169
rect 1223 135 1236 169
rect 1178 119 1236 135
rect 1266 203 1316 267
rect 2036 210 2093 242
rect 2036 204 2048 210
rect 1266 175 1520 203
rect 1266 141 1341 175
rect 1375 141 1475 175
rect 1509 141 1520 175
rect 1266 119 1520 141
rect 1550 119 1598 203
rect 1628 165 1706 203
rect 1628 131 1650 165
rect 1684 131 1706 165
rect 1628 119 1706 131
rect 1736 119 1784 203
rect 1814 170 1871 203
rect 1814 136 1825 170
rect 1859 136 1871 170
rect 1814 119 1871 136
rect 1934 166 1991 204
rect 1934 132 1946 166
rect 1980 132 1991 166
rect 1055 90 1067 119
rect 1009 78 1067 90
rect 1934 94 1991 132
rect 2021 176 2048 204
rect 2082 176 2093 210
rect 2021 138 2093 176
rect 2021 104 2048 138
rect 2082 104 2093 138
rect 2021 94 2093 104
rect 2123 214 2181 242
rect 2123 180 2134 214
rect 2168 180 2181 214
rect 2123 138 2181 180
rect 2123 104 2134 138
rect 2168 104 2181 138
rect 2123 94 2181 104
<< pdiff >>
rect 27 567 85 592
rect 27 533 38 567
rect 72 533 85 567
rect 27 508 85 533
rect 115 567 175 592
rect 115 533 128 567
rect 162 533 175 567
rect 115 508 175 533
rect 205 554 261 592
rect 205 520 219 554
rect 253 547 261 554
rect 1106 580 1161 592
rect 253 520 276 547
rect 205 508 276 520
rect 223 347 276 508
rect 306 398 364 547
rect 306 364 319 398
rect 353 364 364 398
rect 306 347 364 364
rect 418 538 477 547
rect 418 504 430 538
rect 464 504 477 538
rect 418 347 477 504
rect 507 429 584 547
rect 638 527 697 547
rect 638 493 650 527
rect 684 493 697 527
rect 638 463 697 493
rect 727 527 787 547
rect 727 493 740 527
rect 774 493 787 527
rect 727 463 787 493
rect 817 463 865 547
rect 895 527 964 547
rect 895 493 908 527
rect 942 493 964 527
rect 895 463 964 493
rect 994 527 1052 547
rect 994 493 1010 527
rect 1044 493 1052 527
rect 994 463 1052 493
rect 1106 546 1114 580
rect 1148 546 1161 580
rect 1106 506 1161 546
rect 1106 472 1114 506
rect 1148 472 1161 506
rect 507 398 593 429
rect 507 364 551 398
rect 585 364 593 398
rect 507 347 593 364
rect 1106 392 1161 472
rect 1191 580 1347 592
rect 1191 546 1205 580
rect 1239 546 1299 580
rect 1333 546 1347 580
rect 1191 512 1347 546
rect 1191 478 1205 512
rect 1239 478 1299 512
rect 1333 478 1347 512
rect 1191 444 1347 478
rect 1191 410 1205 444
rect 1239 410 1299 444
rect 1333 410 1347 444
rect 1191 392 1347 410
rect 1377 557 1517 592
rect 1377 523 1390 557
rect 1424 523 1470 557
rect 1504 523 1517 557
rect 1377 508 1517 523
rect 1547 508 1601 592
rect 1631 567 1709 592
rect 1631 533 1644 567
rect 1678 533 1709 567
rect 1631 508 1709 533
rect 1739 567 1799 592
rect 1739 533 1752 567
rect 1786 533 1799 567
rect 1739 508 1799 533
rect 1829 567 1884 592
rect 1829 533 1842 567
rect 1876 533 1884 567
rect 1829 508 1884 533
rect 1938 580 1993 592
rect 1938 546 1946 580
rect 1980 546 1993 580
rect 1377 392 1430 508
rect 1938 471 1993 546
rect 1938 437 1946 471
rect 1980 437 1993 471
rect 1938 424 1993 437
rect 2023 580 2094 592
rect 2023 546 2046 580
rect 2080 546 2094 580
rect 2023 470 2094 546
rect 2023 436 2046 470
rect 2080 436 2094 470
rect 2023 424 2094 436
rect 2041 368 2094 424
rect 2124 580 2181 592
rect 2124 546 2137 580
rect 2171 546 2181 580
rect 2124 497 2181 546
rect 2124 463 2137 497
rect 2171 463 2181 497
rect 2124 414 2181 463
rect 2124 380 2137 414
rect 2171 380 2181 414
rect 2124 368 2181 380
<< ndiffc >>
rect 45 97 79 131
rect 225 99 259 133
rect 311 168 345 202
rect 311 86 345 120
rect 535 181 569 215
rect 639 154 673 188
rect 775 154 809 188
rect 417 43 451 77
rect 1021 90 1055 124
rect 1189 210 1223 244
rect 1189 135 1223 169
rect 1341 141 1375 175
rect 1475 141 1509 175
rect 1650 131 1684 165
rect 1825 136 1859 170
rect 1946 132 1980 166
rect 2048 176 2082 210
rect 2048 104 2082 138
rect 2134 180 2168 214
rect 2134 104 2168 138
<< pdiffc >>
rect 38 533 72 567
rect 128 533 162 567
rect 219 520 253 554
rect 319 364 353 398
rect 430 504 464 538
rect 650 493 684 527
rect 740 493 774 527
rect 908 493 942 527
rect 1010 493 1044 527
rect 1114 546 1148 580
rect 1114 472 1148 506
rect 551 364 585 398
rect 1205 546 1239 580
rect 1299 546 1333 580
rect 1205 478 1239 512
rect 1299 478 1333 512
rect 1205 410 1239 444
rect 1299 410 1333 444
rect 1390 523 1424 557
rect 1470 523 1504 557
rect 1644 533 1678 567
rect 1752 533 1786 567
rect 1842 533 1876 567
rect 1946 546 1980 580
rect 1946 437 1980 471
rect 2046 546 2080 580
rect 2046 436 2080 470
rect 2137 546 2171 580
rect 2137 463 2171 497
rect 2137 380 2171 414
<< poly >>
rect 85 592 115 618
rect 175 615 994 645
rect 175 592 205 615
rect 276 547 306 573
rect 477 547 507 573
rect 697 547 727 573
rect 787 547 817 573
rect 865 547 895 573
rect 964 547 994 615
rect 1161 592 1191 618
rect 1347 592 1377 618
rect 1517 592 1547 618
rect 1601 592 1631 618
rect 1709 592 1739 618
rect 1799 592 1829 618
rect 1993 592 2023 618
rect 2094 592 2124 618
rect 85 493 115 508
rect 82 414 118 493
rect 175 448 205 508
rect 57 384 118 414
rect 57 326 87 384
rect 172 332 208 448
rect 697 448 727 463
rect 787 448 817 463
rect 608 418 727 448
rect 769 418 817 448
rect 865 448 895 463
rect 964 448 994 463
rect 276 332 306 347
rect 477 332 507 347
rect 608 332 638 418
rect 769 376 799 418
rect 865 376 922 448
rect 21 310 87 326
rect 21 276 37 310
rect 71 276 87 310
rect 21 242 87 276
rect 21 208 37 242
rect 71 222 87 242
rect 162 299 228 332
rect 162 265 178 299
rect 212 265 228 299
rect 162 237 228 265
rect 270 299 341 332
rect 270 265 291 299
rect 325 265 341 299
rect 270 237 341 265
rect 383 299 638 332
rect 680 360 799 376
rect 680 326 696 360
rect 730 326 799 360
rect 680 310 799 326
rect 841 339 922 376
rect 383 265 399 299
rect 433 265 638 299
rect 383 242 638 265
rect 744 258 774 310
rect 841 305 857 339
rect 891 305 922 339
rect 841 288 922 305
rect 71 208 120 222
rect 21 192 120 208
rect 90 158 120 192
rect 168 158 198 237
rect 270 222 300 237
rect 480 227 510 242
rect 684 228 774 258
rect 684 211 714 228
rect 820 211 850 237
rect 892 211 922 288
rect 964 360 1011 448
rect 1517 493 1547 508
rect 1601 493 1631 508
rect 1709 493 1739 508
rect 1799 493 1829 508
rect 1514 473 1547 493
rect 1462 457 1544 473
rect 1462 423 1478 457
rect 1512 423 1544 457
rect 1161 377 1191 392
rect 1347 377 1377 392
rect 1462 389 1544 423
rect 1158 360 1194 377
rect 964 344 1033 360
rect 964 310 983 344
rect 1017 310 1033 344
rect 964 294 1033 310
rect 1075 344 1194 360
rect 1075 310 1091 344
rect 1125 310 1194 344
rect 1075 294 1194 310
rect 1236 344 1302 360
rect 1236 310 1252 344
rect 1286 310 1302 344
rect 1236 294 1302 310
rect 964 226 1011 294
rect 1148 267 1178 294
rect 1236 267 1266 294
rect 1344 291 1380 377
rect 1462 355 1478 389
rect 1512 355 1544 389
rect 1462 339 1544 355
rect 1598 467 1634 493
rect 1598 451 1664 467
rect 1598 417 1614 451
rect 1648 417 1664 451
rect 1598 401 1664 417
rect 1344 275 1484 291
rect 964 211 994 226
rect 684 101 714 127
rect 90 48 120 74
rect 168 48 198 74
rect 270 48 300 74
rect 480 51 510 79
rect 820 51 850 127
rect 892 101 922 127
rect 964 101 994 127
rect 1344 261 1366 275
rect 1350 241 1366 261
rect 1400 241 1434 275
rect 1468 255 1484 275
rect 1468 241 1550 255
rect 1350 225 1550 241
rect 1520 203 1550 225
rect 1598 203 1628 401
rect 1706 359 1742 493
rect 1796 409 1832 493
rect 1993 409 2023 424
rect 1796 379 2026 409
rect 1796 359 1850 379
rect 1676 343 1742 359
rect 1676 309 1692 343
rect 1726 309 1742 343
rect 1676 293 1742 309
rect 1784 343 1850 359
rect 2094 353 2124 368
rect 1784 309 1800 343
rect 1834 309 1850 343
rect 2091 330 2127 353
rect 1706 203 1736 293
rect 1784 275 1850 309
rect 1784 241 1800 275
rect 1834 255 1850 275
rect 2063 314 2129 330
rect 2063 280 2079 314
rect 2113 280 2129 314
rect 2063 264 2129 280
rect 1834 241 2021 255
rect 2093 242 2123 264
rect 1784 225 2021 241
rect 1784 203 1814 225
rect 1991 204 2021 225
rect 1148 93 1178 119
rect 1236 51 1266 119
rect 1520 93 1550 119
rect 1598 93 1628 119
rect 1706 93 1736 119
rect 1784 93 1814 119
rect 1991 68 2021 94
rect 2093 68 2123 94
rect 480 21 1266 51
<< polycont >>
rect 37 276 71 310
rect 37 208 71 242
rect 178 265 212 299
rect 291 265 325 299
rect 696 326 730 360
rect 399 265 433 299
rect 857 305 891 339
rect 1478 423 1512 457
rect 983 310 1017 344
rect 1091 310 1125 344
rect 1252 310 1286 344
rect 1478 355 1512 389
rect 1614 417 1648 451
rect 1366 241 1400 275
rect 1434 241 1468 275
rect 1692 309 1726 343
rect 1800 309 1834 343
rect 1800 241 1834 275
rect 2079 280 2113 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 22 567 88 649
rect 22 533 38 567
rect 72 533 88 567
rect 22 504 88 533
rect 128 567 174 596
rect 162 533 174 567
rect 128 470 174 533
rect 208 554 274 649
rect 208 520 219 554
rect 253 520 274 554
rect 208 504 274 520
rect 414 538 480 649
rect 414 504 430 538
rect 464 504 480 538
rect 634 527 684 547
rect 634 493 650 527
rect 634 470 684 493
rect 108 436 684 470
rect 724 527 815 547
rect 724 493 740 527
rect 774 493 815 527
rect 724 436 815 493
rect 892 527 958 649
rect 1098 580 1164 649
rect 892 493 908 527
rect 942 493 958 527
rect 892 462 958 493
rect 994 527 1060 547
rect 994 493 1010 527
rect 1044 493 1060 527
rect 21 310 74 430
rect 21 276 37 310
rect 71 276 74 310
rect 21 242 74 276
rect 21 208 37 242
rect 71 208 74 242
rect 21 192 74 208
rect 108 158 142 436
rect 303 398 433 402
rect 303 364 319 398
rect 353 364 433 398
rect 176 350 257 356
rect 176 316 223 350
rect 176 299 257 316
rect 176 265 178 299
rect 212 265 257 299
rect 176 249 257 265
rect 291 299 353 330
rect 325 265 353 299
rect 291 236 353 265
rect 387 299 433 364
rect 387 265 399 299
rect 387 202 433 265
rect 295 168 311 202
rect 345 168 433 202
rect 29 131 142 158
rect 29 97 45 131
rect 79 97 142 131
rect 29 70 142 97
rect 209 133 259 162
rect 209 99 225 133
rect 209 17 259 99
rect 295 133 433 168
rect 467 145 501 436
rect 775 428 815 436
rect 994 428 1060 493
rect 1098 546 1114 580
rect 1148 546 1164 580
rect 1098 506 1164 546
rect 1098 472 1114 506
rect 1148 472 1164 506
rect 1198 580 1340 596
rect 1198 546 1205 580
rect 1239 546 1299 580
rect 1333 546 1340 580
rect 1198 512 1340 546
rect 1198 478 1205 512
rect 1239 478 1299 512
rect 1333 478 1340 512
rect 1374 557 1520 573
rect 1374 523 1390 557
rect 1424 523 1470 557
rect 1504 541 1520 557
rect 1628 567 1694 649
rect 1504 523 1580 541
rect 1374 507 1580 523
rect 1198 444 1340 478
rect 1198 428 1205 444
rect 535 398 741 402
rect 535 364 551 398
rect 585 364 741 398
rect 535 360 741 364
rect 535 326 696 360
rect 730 326 741 360
rect 535 249 741 326
rect 535 215 588 249
rect 569 181 588 215
rect 535 165 588 181
rect 623 188 673 215
rect 623 154 639 188
rect 467 141 507 145
rect 467 137 510 141
rect 295 120 361 133
rect 467 131 515 137
rect 623 131 673 154
rect 467 125 673 131
rect 471 121 673 125
rect 295 86 311 120
rect 345 86 361 120
rect 474 119 673 121
rect 479 113 673 119
rect 482 109 673 113
rect 483 105 673 109
rect 488 97 673 105
rect 707 93 741 249
rect 775 394 1139 428
rect 775 188 815 394
rect 855 339 931 355
rect 855 305 857 339
rect 891 305 931 339
rect 855 260 931 305
rect 971 350 1031 360
rect 971 344 991 350
rect 971 310 983 344
rect 1025 316 1031 350
rect 1017 310 1031 316
rect 971 294 1031 310
rect 1067 344 1139 394
rect 1067 310 1091 344
rect 1125 310 1139 344
rect 1067 294 1139 310
rect 1173 410 1205 428
rect 1239 410 1299 444
rect 1333 410 1340 444
rect 1173 394 1340 410
rect 1462 457 1512 473
rect 1462 423 1478 457
rect 1173 260 1207 394
rect 1462 389 1512 423
rect 1462 360 1478 389
rect 1241 355 1478 360
rect 1241 344 1512 355
rect 1241 310 1252 344
rect 1286 326 1512 344
rect 1286 310 1302 326
rect 1241 294 1302 310
rect 1350 275 1484 291
rect 855 244 1239 260
rect 1350 259 1366 275
rect 855 226 1189 244
rect 1173 210 1189 226
rect 1223 210 1239 244
rect 809 154 815 188
rect 775 127 815 154
rect 937 158 1139 192
rect 937 93 971 158
rect 295 70 361 86
rect 404 77 451 93
rect 404 43 417 77
rect 707 51 971 93
rect 1005 90 1021 124
rect 1055 90 1071 124
rect 404 17 451 43
rect 1005 17 1071 90
rect 1105 85 1139 158
rect 1173 169 1239 210
rect 1173 135 1189 169
rect 1223 135 1239 169
rect 1173 119 1239 135
rect 1273 241 1366 259
rect 1400 241 1434 275
rect 1468 241 1484 275
rect 1273 225 1484 241
rect 1546 259 1580 507
rect 1628 533 1644 567
rect 1678 533 1694 567
rect 1628 504 1694 533
rect 1736 567 1802 596
rect 1736 533 1752 567
rect 1786 533 1802 567
rect 1736 467 1802 533
rect 1842 567 1892 649
rect 1876 533 1892 567
rect 1842 504 1892 533
rect 1930 580 1996 596
rect 1930 546 1946 580
rect 1980 546 1996 580
rect 1930 471 1996 546
rect 1614 451 1810 467
rect 1930 461 1946 471
rect 1648 427 1810 451
rect 1980 437 1996 471
rect 1648 417 1912 427
rect 1614 393 1912 417
rect 1657 350 1742 359
rect 1657 316 1663 350
rect 1697 343 1742 350
rect 1657 309 1692 316
rect 1726 309 1742 343
rect 1657 293 1742 309
rect 1784 343 1844 359
rect 1784 309 1800 343
rect 1834 309 1844 343
rect 1784 275 1844 309
rect 1784 259 1800 275
rect 1546 241 1800 259
rect 1834 241 1844 275
rect 1546 225 1844 241
rect 1273 85 1307 225
rect 1546 191 1580 225
rect 1878 191 1912 393
rect 1341 175 1580 191
rect 1375 141 1475 175
rect 1509 141 1580 175
rect 1341 125 1580 141
rect 1623 165 1711 181
rect 1623 131 1650 165
rect 1684 131 1711 165
rect 1105 51 1307 85
rect 1623 17 1711 131
rect 1809 170 1912 191
rect 1809 136 1825 170
rect 1859 136 1912 170
rect 1809 115 1912 136
rect 1946 330 1996 437
rect 2030 580 2080 649
rect 2030 546 2046 580
rect 2030 470 2080 546
rect 2030 436 2046 470
rect 2030 420 2080 436
rect 2121 580 2191 596
rect 2121 546 2137 580
rect 2171 546 2191 580
rect 2121 497 2191 546
rect 2121 463 2137 497
rect 2171 463 2191 497
rect 2121 414 2191 463
rect 2121 380 2137 414
rect 2171 380 2191 414
rect 2121 364 2191 380
rect 1946 314 2123 330
rect 1946 280 2079 314
rect 2113 280 2123 314
rect 1946 264 2123 280
rect 1946 166 1996 264
rect 2157 230 2191 364
rect 1980 132 1996 166
rect 1946 106 1996 132
rect 2032 210 2082 226
rect 2032 176 2048 210
rect 2032 138 2082 176
rect 2032 104 2048 138
rect 2032 17 2082 104
rect 2118 214 2191 230
rect 2118 180 2134 214
rect 2168 180 2191 214
rect 2118 138 2191 180
rect 2118 104 2134 138
rect 2168 104 2191 138
rect 2118 88 2191 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 316 257 350
rect 991 344 1025 350
rect 991 316 1017 344
rect 1017 316 1025 344
rect 1663 343 1697 350
rect 1663 316 1692 343
rect 1692 316 1697 343
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 979 350 1037 356
rect 979 347 991 350
rect 257 319 991 347
rect 257 316 269 319
rect 211 310 269 316
rect 979 316 991 319
rect 1025 347 1037 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1025 319 1663 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel comment s 566 630 566 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrtn_1
flabel comment s 619 296 619 296 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 223 316 257 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew
flabel corelocali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew
flabel corelocali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 8 nsew
flabel corelocali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew
flabel corelocali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 666
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 2585946
string GDS_START 2569258
<< end >>
