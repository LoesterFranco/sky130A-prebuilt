magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 736 561
rect 18 298 77 527
rect 18 17 77 181
rect 111 127 157 467
rect 200 366 251 527
rect 391 438 446 527
rect 296 209 362 255
rect 396 209 490 255
rect 524 209 614 255
rect 652 209 719 255
rect 111 51 155 127
rect 189 17 359 89
rect 562 17 617 105
rect 0 -17 736 17
<< obsli1 >>
rect 291 404 357 493
rect 493 404 559 493
rect 291 368 559 404
rect 651 332 717 465
rect 200 298 717 332
rect 200 175 262 298
rect 200 139 717 175
rect 455 55 521 139
rect 651 55 717 139
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 396 209 490 255 6 A1
port 1 nsew signal input
rlabel locali s 296 209 362 255 6 A2
port 2 nsew signal input
rlabel locali s 524 209 614 255 6 B1
port 3 nsew signal input
rlabel locali s 652 209 719 255 6 C1
port 4 nsew signal input
rlabel locali s 111 127 157 467 6 X
port 5 nsew signal output
rlabel locali s 111 51 155 127 6 X
port 5 nsew signal output
rlabel locali s 562 17 617 105 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 189 17 359 89 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 18 17 77 181 6 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 0 -17 736 17 8 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel locali s 391 438 446 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 200 366 251 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 18 298 77 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3925878
string GDS_START 3919314
<< end >>
