magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 465 47 495 177
rect 663 47 693 177
rect 757 47 787 177
rect 849 47 879 177
rect 944 47 974 177
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 655 297 691 497
rect 749 297 785 497
rect 851 297 887 497
rect 946 297 982 497
<< ndiff >>
rect 27 119 89 177
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 177
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 165 277 177
rect 213 131 223 165
rect 257 131 277 165
rect 213 47 277 131
rect 307 161 371 177
rect 307 127 317 161
rect 351 127 371 161
rect 307 93 371 127
rect 307 59 317 93
rect 351 59 371 93
rect 307 47 371 59
rect 401 109 465 177
rect 401 75 411 109
rect 445 75 465 109
rect 401 47 465 75
rect 495 93 547 177
rect 495 59 505 93
rect 539 59 547 93
rect 495 47 547 59
rect 601 93 663 177
rect 601 59 609 93
rect 643 59 663 93
rect 601 47 663 59
rect 693 165 757 177
rect 693 131 703 165
rect 737 131 757 165
rect 693 47 757 131
rect 787 93 849 177
rect 787 59 797 93
rect 831 59 849 93
rect 787 47 849 59
rect 879 165 944 177
rect 879 131 899 165
rect 933 131 944 165
rect 879 47 944 131
rect 974 93 1075 177
rect 974 59 1033 93
rect 1067 59 1075 93
rect 974 47 1075 59
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 297 81 443
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 297 175 451
rect 211 401 269 497
rect 211 367 223 401
rect 257 367 269 401
rect 211 297 269 367
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 297 363 451
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 297 457 443
rect 493 485 547 497
rect 493 451 505 485
rect 539 451 547 485
rect 493 297 547 451
rect 601 485 655 497
rect 601 451 609 485
rect 643 451 655 485
rect 601 297 655 451
rect 691 343 749 497
rect 691 309 703 343
rect 737 309 749 343
rect 691 297 749 309
rect 785 485 851 497
rect 785 451 801 485
rect 835 451 851 485
rect 785 297 851 451
rect 887 417 946 497
rect 887 383 900 417
rect 934 383 946 417
rect 887 297 946 383
rect 982 485 1075 497
rect 982 451 995 485
rect 1029 451 1075 485
rect 982 297 1075 451
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 131 257 165
rect 317 127 351 161
rect 317 59 351 93
rect 411 75 445 109
rect 505 59 539 93
rect 609 59 643 93
rect 703 131 737 165
rect 797 59 831 93
rect 899 131 933 165
rect 1033 59 1067 93
<< pdiffc >>
rect 35 443 69 477
rect 129 451 163 485
rect 223 367 257 401
rect 317 451 351 485
rect 411 443 445 477
rect 505 451 539 485
rect 609 451 643 485
rect 703 309 737 343
rect 801 451 835 485
rect 900 383 934 417
rect 995 451 1029 485
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 655 497 691 523
rect 749 497 785 523
rect 851 497 887 523
rect 946 497 982 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 655 282 691 297
rect 749 282 785 297
rect 851 282 887 297
rect 946 282 982 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 76 249 307 265
rect 76 215 86 249
rect 120 215 307 249
rect 76 199 307 215
rect 358 249 495 265
rect 653 265 693 282
rect 747 265 787 282
rect 849 265 889 282
rect 944 265 984 282
rect 653 259 794 265
rect 358 215 377 249
rect 411 215 495 249
rect 358 205 495 215
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 199
rect 371 177 401 205
rect 465 177 495 205
rect 544 249 794 259
rect 544 215 560 249
rect 594 215 628 249
rect 662 215 706 249
rect 740 215 794 249
rect 544 199 794 215
rect 849 249 1032 265
rect 849 215 973 249
rect 1007 215 1032 249
rect 849 199 1032 215
rect 663 177 693 199
rect 757 177 787 199
rect 849 177 879 199
rect 944 177 974 199
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 465 21 495 47
rect 663 21 693 47
rect 757 21 787 47
rect 849 21 879 47
rect 944 21 974 47
<< polycont >>
rect 86 215 120 249
rect 377 215 411 249
rect 560 215 594 249
rect 628 215 662 249
rect 706 215 740 249
rect 973 215 1007 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 291 485 367 527
rect 291 451 317 485
rect 351 451 367 485
rect 411 477 456 493
rect 17 427 69 443
rect 445 443 456 477
rect 411 427 456 443
rect 505 485 555 527
rect 539 451 555 485
rect 593 451 609 485
rect 643 451 801 485
rect 835 451 995 485
rect 1029 451 1085 485
rect 505 435 555 451
rect 17 333 52 427
rect 422 401 456 427
rect 593 401 900 417
rect 197 367 223 401
rect 257 367 377 401
rect 422 383 900 401
rect 934 383 950 417
rect 422 367 627 383
rect 343 333 377 367
rect 1040 357 1085 451
rect 677 333 703 343
rect 17 299 309 333
rect 343 309 703 333
rect 737 309 753 343
rect 343 299 753 309
rect 17 135 52 299
rect 265 265 309 299
rect 86 249 166 265
rect 120 215 166 249
rect 265 249 437 265
rect 265 231 377 249
rect 361 215 377 231
rect 411 215 437 249
rect 544 249 805 255
rect 544 215 560 249
rect 594 215 628 249
rect 662 215 706 249
rect 740 215 805 249
rect 942 249 1017 323
rect 942 215 973 249
rect 1007 215 1017 249
rect 86 199 166 215
rect 942 199 1017 215
rect 126 145 166 199
rect 223 165 234 187
rect 268 153 271 187
rect 17 119 69 135
rect 17 85 35 119
rect 257 131 271 153
rect 223 115 271 131
rect 317 161 367 177
rect 351 127 367 161
rect 17 69 69 85
rect 103 93 177 109
rect 103 59 129 93
rect 163 59 177 93
rect 103 17 177 59
rect 317 93 367 127
rect 351 59 367 93
rect 411 165 753 181
rect 411 147 703 165
rect 411 109 445 147
rect 677 131 703 147
rect 737 131 753 165
rect 874 165 901 187
rect 874 153 899 165
rect 840 131 899 153
rect 933 131 949 165
rect 411 59 445 75
rect 505 93 539 109
rect 1051 93 1085 357
rect 593 59 609 93
rect 643 59 797 93
rect 831 59 1033 93
rect 1067 59 1085 93
rect 317 17 367 59
rect 505 17 539 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 234 165 268 187
rect 234 153 257 165
rect 257 153 268 165
rect 840 153 874 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 222 187 280 193
rect 222 153 234 187
rect 268 184 280 187
rect 828 187 896 193
rect 828 184 840 187
rect 268 156 840 184
rect 268 153 280 156
rect 222 147 280 153
rect 828 153 840 156
rect 874 153 896 187
rect 828 147 896 153
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel corelocali s 1040 425 1074 459 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 952 289 986 323 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 952 221 986 255 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel corelocali s 1040 357 1074 391 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel corelocali s 669 221 703 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 576 221 610 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 764 221 798 255 0 FreeSans 200 0 0 0 A0
port 1 nsew
flabel corelocali s 132 221 166 255 0 FreeSans 200 0 0 0 S
port 3 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nbase s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
rlabel comment s 0 0 0 0 4 mux2i_2
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 2174066
string GDS_START 2165604
<< end >>
