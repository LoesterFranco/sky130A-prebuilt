magic
tech sky130A
magscale 1 2
timestamp 1604502729
<< locali >>
rect 257 430 323 596
rect 457 430 527 596
rect 257 378 527 430
rect 257 364 655 378
rect 323 344 655 364
rect 89 236 163 310
rect 197 236 263 310
rect 305 236 371 310
rect 409 236 479 310
rect 621 210 655 344
rect 581 70 655 210
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 21 364 116 540
rect 157 364 223 649
rect 357 464 423 649
rect 561 412 627 649
rect 21 202 55 364
rect 513 244 587 310
rect 513 202 547 244
rect 21 168 547 202
rect 21 136 130 168
rect 171 17 237 134
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 89 236 163 310 6 A_N
port 1 nsew signal input
rlabel locali s 409 236 479 310 6 B
port 2 nsew signal input
rlabel locali s 305 236 371 310 6 C
port 3 nsew signal input
rlabel locali s 197 236 263 310 6 D
port 4 nsew signal input
rlabel locali s 621 210 655 344 6 Y
port 5 nsew signal output
rlabel locali s 581 70 655 210 6 Y
port 5 nsew signal output
rlabel locali s 457 430 527 596 6 Y
port 5 nsew signal output
rlabel locali s 323 344 655 364 6 Y
port 5 nsew signal output
rlabel locali s 257 430 323 596 6 Y
port 5 nsew signal output
rlabel locali s 257 378 527 430 6 Y
port 5 nsew signal output
rlabel locali s 257 364 655 378 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1452656
string GDS_START 1446650
<< end >>
