magic
tech sky130A
magscale 1 2
timestamp 1601050082
<< locali >>
rect 121 370 460 420
rect 121 302 284 370
rect 25 101 71 134
rect 25 51 125 101
rect 250 236 284 302
rect 889 290 1040 356
rect 250 202 483 236
rect 250 96 311 202
rect 433 96 483 202
rect 787 51 853 134
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 21 488 87 596
rect 124 522 190 649
rect 304 522 370 649
rect 484 522 550 649
rect 588 581 818 615
rect 21 454 528 488
rect 21 255 87 454
rect 494 404 528 454
rect 588 438 654 581
rect 494 370 658 404
rect 21 168 123 255
rect 159 17 209 255
rect 318 270 551 336
rect 592 290 658 370
rect 517 256 551 270
rect 694 256 744 547
rect 784 424 818 581
rect 858 458 908 649
rect 948 424 1014 596
rect 1054 458 1104 649
rect 1144 424 1194 596
rect 784 390 1194 424
rect 784 388 818 390
rect 1144 388 1194 390
rect 517 222 1007 256
rect 347 17 397 168
rect 519 17 569 188
rect 617 119 683 222
rect 719 17 753 188
rect 887 85 921 188
rect 957 119 1007 222
rect 1043 85 1109 255
rect 887 51 1109 85
rect 1145 17 1195 255
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel locali s 889 290 1040 356 6 A1
port 1 nsew signal input
rlabel locali s 787 51 853 134 6 A2
port 2 nsew signal input
rlabel locali s 25 101 71 134 6 B1_N
port 3 nsew signal input
rlabel locali s 25 51 125 101 6 B1_N
port 3 nsew signal input
rlabel locali s 433 96 483 202 6 X
port 4 nsew signal output
rlabel locali s 250 236 284 302 6 X
port 4 nsew signal output
rlabel locali s 250 202 483 236 6 X
port 4 nsew signal output
rlabel locali s 250 96 311 202 6 X
port 4 nsew signal output
rlabel locali s 121 370 460 420 6 X
port 4 nsew signal output
rlabel locali s 121 302 284 370 6 X
port 4 nsew signal output
rlabel metal1 s 0 -49 1248 49 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 617 1248 715 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string GDS_END 4042894
string GDS_START 4032920
<< end >>
