magic
tech sky130A
magscale 1 2
timestamp 1599588220
<< locali >>
rect 0 527 1656 561
rect 17 288 73 493
rect 107 443 174 527
rect 645 447 711 527
rect 1479 455 1546 527
rect 17 185 66 288
rect 17 70 69 185
rect 103 17 153 105
rect 323 215 436 265
rect 695 17 729 173
rect 1245 289 1361 323
rect 1245 199 1279 289
rect 1409 215 1491 265
rect 1495 17 1529 113
rect 0 -17 1656 17
<< obsli1 >>
rect 210 447 504 481
rect 778 455 1397 489
rect 210 409 244 447
rect 778 413 812 455
rect 107 375 244 409
rect 312 379 812 413
rect 107 265 141 375
rect 187 307 504 341
rect 100 199 141 265
rect 106 173 141 199
rect 106 139 221 173
rect 187 85 221 139
rect 255 119 289 307
rect 470 265 504 307
rect 538 323 615 339
rect 538 305 581 323
rect 559 289 581 305
rect 559 275 615 289
rect 470 199 525 265
rect 349 159 425 181
rect 559 159 593 275
rect 649 241 683 379
rect 729 289 813 343
rect 349 125 593 159
rect 627 207 683 241
rect 627 91 661 207
rect 765 187 813 289
rect 414 85 501 91
rect 187 51 501 85
rect 535 57 661 91
rect 799 153 813 187
rect 765 83 813 153
rect 849 119 883 421
rect 917 178 951 455
rect 1580 421 1639 493
rect 987 323 1070 409
rect 1177 387 1639 421
rect 987 289 1041 323
rect 1075 289 1143 323
rect 990 199 1075 254
rect 1033 187 1075 199
rect 917 165 959 178
rect 917 144 999 165
rect 925 131 999 144
rect 849 85 857 119
rect 891 85 931 97
rect 849 53 931 85
rect 965 64 999 131
rect 1033 153 1041 187
rect 1033 126 1075 153
rect 1109 85 1143 289
rect 1177 119 1211 387
rect 1542 375 1639 387
rect 1395 299 1559 341
rect 1525 265 1559 299
rect 1313 189 1375 255
rect 1525 199 1571 265
rect 1313 187 1354 189
rect 1313 153 1317 187
rect 1351 153 1354 187
rect 1525 181 1559 199
rect 1313 146 1354 153
rect 1411 150 1559 181
rect 1403 147 1559 150
rect 1403 119 1461 147
rect 1245 85 1338 93
rect 1109 51 1338 85
rect 1403 85 1409 119
rect 1443 85 1461 119
rect 1605 117 1639 375
rect 1403 59 1461 85
rect 1579 51 1639 117
<< obsli1c >>
rect 581 289 615 323
rect 765 153 799 187
rect 1041 289 1075 323
rect 857 85 891 119
rect 1041 153 1075 187
rect 1317 153 1351 187
rect 1409 85 1443 119
<< metal1 >>
rect 0 496 1656 592
rect 0 -48 1656 48
<< obsm1 >>
rect 569 323 627 329
rect 569 289 581 323
rect 615 320 627 323
rect 1029 323 1087 329
rect 1029 320 1041 323
rect 615 292 1041 320
rect 615 289 627 292
rect 569 283 627 289
rect 1029 289 1041 292
rect 1075 289 1087 323
rect 1029 283 1087 289
rect 753 187 811 193
rect 753 153 765 187
rect 799 184 811 187
rect 1029 187 1087 193
rect 1029 184 1041 187
rect 799 156 1041 184
rect 799 153 811 156
rect 753 147 811 153
rect 1029 153 1041 156
rect 1075 184 1087 187
rect 1305 187 1363 193
rect 1305 184 1317 187
rect 1075 156 1317 184
rect 1075 153 1087 156
rect 1029 147 1087 153
rect 1305 153 1317 156
rect 1351 153 1363 187
rect 1305 147 1363 153
rect 845 119 903 125
rect 845 85 857 119
rect 891 116 903 119
rect 1397 119 1455 125
rect 1397 116 1409 119
rect 891 88 1409 116
rect 891 85 903 88
rect 845 79 903 85
rect 1397 85 1409 88
rect 1443 85 1455 119
rect 1397 79 1455 85
<< labels >>
rlabel locali s 1409 215 1491 265 6 A
port 1 nsew signal input
rlabel locali s 1245 289 1361 323 6 B
port 2 nsew signal input
rlabel locali s 1245 199 1279 289 6 B
port 2 nsew signal input
rlabel locali s 323 215 436 265 6 C
port 3 nsew signal input
rlabel locali s 17 288 73 493 6 X
port 4 nsew signal output
rlabel locali s 17 185 66 288 6 X
port 4 nsew signal output
rlabel locali s 17 70 69 185 6 X
port 4 nsew signal output
rlabel locali s 1495 17 1529 113 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 695 17 729 173 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 153 105 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1656 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1656 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1479 455 1546 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 645 447 711 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 107 443 174 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1656 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 496 1656 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 604160
string GDS_START 592554
<< end >>
