magic
tech sky130A
magscale 1 2
timestamp 1601050043
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 84 -17 128 17
<< scnmos >>
rect 79 47 109 151
rect 215 47 245 131
rect 317 47 347 131
rect 448 47 478 131
rect 649 47 679 131
rect 773 47 803 151
<< pmoshvt >>
rect 81 297 117 497
rect 207 309 243 497
rect 326 309 362 497
rect 563 309 599 497
rect 651 309 687 497
rect 765 309 801 497
<< ndiff >>
rect 27 112 79 151
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 109 131 171 151
rect 723 131 773 151
rect 109 93 215 131
rect 109 59 129 93
rect 163 59 215 93
rect 109 47 215 59
rect 245 47 317 131
rect 347 108 448 131
rect 347 74 357 108
rect 391 74 448 108
rect 347 47 448 74
rect 478 47 649 131
rect 679 89 773 131
rect 679 55 709 89
rect 743 55 773 89
rect 679 47 773 55
rect 803 108 855 151
rect 803 74 813 108
rect 847 74 855 108
rect 803 47 855 74
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 207 497
rect 117 451 129 485
rect 163 451 207 485
rect 117 417 207 451
rect 117 383 129 417
rect 163 383 207 417
rect 117 349 207 383
rect 117 315 129 349
rect 163 315 207 349
rect 117 309 207 315
rect 243 309 326 497
rect 362 425 563 497
rect 362 391 374 425
rect 408 391 449 425
rect 483 391 517 425
rect 551 391 563 425
rect 362 309 563 391
rect 599 309 651 497
rect 687 485 765 497
rect 687 451 717 485
rect 751 451 765 485
rect 687 417 765 451
rect 687 383 717 417
rect 751 383 765 417
rect 687 309 765 383
rect 801 485 859 497
rect 801 451 813 485
rect 847 451 859 485
rect 801 417 859 451
rect 801 383 813 417
rect 847 383 859 417
rect 801 309 859 383
rect 117 297 171 309
<< ndiffc >>
rect 35 78 69 112
rect 129 59 163 93
rect 357 74 391 108
rect 709 55 743 89
rect 813 74 847 108
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 374 391 408 425
rect 449 391 483 425
rect 517 391 551 425
rect 717 451 751 485
rect 717 383 751 417
rect 813 451 847 485
rect 813 383 847 417
<< poly >>
rect 81 497 117 523
rect 207 497 243 523
rect 326 497 362 523
rect 563 497 599 523
rect 651 497 687 523
rect 765 497 801 523
rect 81 282 117 297
rect 207 294 243 309
rect 326 294 362 309
rect 563 294 599 309
rect 651 294 687 309
rect 765 294 801 309
rect 79 265 119 282
rect 205 265 245 294
rect 79 249 147 265
rect 79 215 103 249
rect 137 215 147 249
rect 79 199 147 215
rect 189 249 245 265
rect 324 264 488 294
rect 561 277 601 294
rect 189 215 199 249
rect 233 215 245 249
rect 448 229 488 264
rect 547 261 601 277
rect 189 199 245 215
rect 79 151 109 199
rect 215 131 245 199
rect 317 212 406 222
rect 317 178 356 212
rect 390 178 406 212
rect 317 168 406 178
rect 448 213 502 229
rect 448 179 458 213
rect 492 179 502 213
rect 547 227 557 261
rect 591 227 601 261
rect 547 211 601 227
rect 649 237 689 294
rect 763 277 803 294
rect 751 261 805 277
rect 649 221 709 237
rect 317 131 347 168
rect 448 163 502 179
rect 649 187 665 221
rect 699 187 709 221
rect 751 227 761 261
rect 795 227 805 261
rect 751 211 805 227
rect 649 171 709 187
rect 448 131 478 163
rect 649 131 679 171
rect 773 151 803 211
rect 79 21 109 47
rect 215 21 245 47
rect 317 21 347 47
rect 448 21 478 47
rect 649 21 679 47
rect 773 21 803 47
<< polycont >>
rect 103 215 137 249
rect 199 215 233 249
rect 356 178 390 212
rect 458 179 492 213
rect 557 227 591 261
rect 665 187 699 221
rect 761 227 795 261
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 485 85 493
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 18 315 35 349
rect 69 315 85 349
rect 18 299 85 315
rect 129 485 163 527
rect 129 417 163 451
rect 129 349 163 383
rect 129 299 163 315
rect 214 459 683 493
rect 18 112 69 299
rect 214 265 254 459
rect 103 249 137 265
rect 103 165 137 215
rect 199 249 254 265
rect 233 215 254 249
rect 199 199 254 215
rect 288 391 374 425
rect 408 391 449 425
rect 483 391 517 425
rect 551 391 577 425
rect 288 165 322 391
rect 103 131 322 165
rect 356 323 615 357
rect 356 212 390 323
rect 356 162 390 178
rect 458 213 523 283
rect 492 179 523 213
rect 18 78 35 112
rect 287 124 322 131
rect 287 108 391 124
rect 18 51 69 78
rect 103 93 179 97
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 287 74 357 108
rect 287 51 391 74
rect 458 51 523 179
rect 557 261 615 323
rect 649 326 683 459
rect 717 485 763 527
rect 751 451 763 485
rect 717 417 763 451
rect 751 383 763 417
rect 717 367 763 383
rect 797 485 877 493
rect 797 451 813 485
rect 847 451 877 485
rect 797 417 877 451
rect 797 383 813 417
rect 847 383 877 417
rect 797 367 877 383
rect 649 288 799 326
rect 591 227 615 261
rect 761 261 799 288
rect 557 51 615 227
rect 665 221 699 237
rect 795 227 799 261
rect 761 211 799 227
rect 665 173 699 187
rect 843 173 877 367
rect 665 139 877 173
rect 807 108 856 139
rect 650 89 753 105
rect 650 55 709 89
rect 743 55 753 89
rect 650 17 753 55
rect 807 74 813 108
rect 847 74 856 108
rect 807 51 856 74
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel corelocali s 672 289 706 323 0 FreeSans 250 0 0 0 S
port 3 nsew
flabel corelocali s 581 153 615 187 0 FreeSans 250 0 0 0 A1
port 2 nsew
flabel corelocali s 581 221 615 255 0 FreeSans 250 0 0 0 A1
port 2 nsew
flabel corelocali s 489 221 523 255 0 FreeSans 250 0 0 0 A0
port 1 nsew
flabel corelocali s 30 85 64 119 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 30 357 64 391 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 30 425 64 459 0 FreeSans 250 0 0 0 X
port 8 nsew
flabel corelocali s 761 289 795 323 0 FreeSans 250 0 0 0 S
port 3 nsew
flabel nbase s 74 527 108 561 0 FreeSans 250 0 0 0 VPB
port 6 nsew
flabel pwell s 84 -17 128 17 0 FreeSans 250 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 clkmux2_1
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3276240
string GDS_START 3269040
<< end >>
