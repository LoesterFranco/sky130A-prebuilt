magic
tech sky130A
magscale 1 2
timestamp 1604502697
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 89 47 119 131
rect 173 47 203 131
rect 277 47 307 131
rect 361 47 391 131
rect 464 47 494 131
rect 549 47 579 131
rect 653 47 683 131
rect 737 47 767 131
<< pmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
<< ndiff >>
rect 27 93 89 131
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 106 173 131
rect 119 72 129 106
rect 163 72 173 106
rect 119 47 173 72
rect 203 106 277 131
rect 203 72 223 106
rect 257 72 277 106
rect 203 47 277 72
rect 307 106 361 131
rect 307 72 317 106
rect 351 72 361 106
rect 307 47 361 72
rect 391 97 464 131
rect 391 63 411 97
rect 445 63 464 97
rect 391 47 464 63
rect 494 106 549 131
rect 494 72 505 106
rect 539 72 549 106
rect 494 47 549 72
rect 579 97 653 131
rect 579 63 599 97
rect 633 63 653 97
rect 579 47 653 63
rect 683 106 737 131
rect 683 72 693 106
rect 727 72 737 106
rect 683 47 737 72
rect 767 97 829 131
rect 767 63 787 97
rect 821 63 829 97
rect 767 47 829 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 349 269 383
rect 211 315 223 349
rect 257 315 269 349
rect 211 297 269 315
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 829 497
rect 775 451 787 485
rect 821 451 829 485
rect 775 417 829 451
rect 775 383 787 417
rect 821 383 829 417
rect 775 297 829 383
<< ndiffc >>
rect 35 59 69 93
rect 129 72 163 106
rect 223 72 257 106
rect 317 72 351 106
rect 411 63 445 97
rect 505 72 539 106
rect 599 63 633 97
rect 693 72 727 106
rect 787 63 821 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 223 315 257 349
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 787 383 821 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 79 265 119 282
rect 173 265 213 282
rect 21 249 213 265
rect 21 215 37 249
rect 71 215 213 249
rect 21 199 213 215
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 267 249 777 265
rect 267 215 288 249
rect 322 215 356 249
rect 390 215 424 249
rect 458 215 492 249
rect 526 215 560 249
rect 594 215 628 249
rect 662 215 777 249
rect 267 199 777 215
rect 89 131 119 199
rect 173 131 203 199
rect 277 131 307 199
rect 361 131 391 199
rect 464 131 494 199
rect 549 131 579 199
rect 653 131 683 199
rect 737 131 767 199
rect 89 21 119 47
rect 173 21 203 47
rect 277 21 307 47
rect 361 21 391 47
rect 464 21 494 47
rect 549 21 579 47
rect 653 21 683 47
rect 737 21 767 47
<< polycont >>
rect 37 215 71 249
rect 288 215 322 249
rect 356 215 390 249
rect 424 215 458 249
rect 492 215 526 249
rect 560 215 594 249
rect 628 215 662 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 19 485 79 527
rect 19 451 35 485
rect 69 451 79 485
rect 19 417 79 451
rect 19 383 35 417
rect 69 383 79 417
rect 19 349 79 383
rect 19 315 35 349
rect 69 315 79 349
rect 19 299 79 315
rect 113 485 179 493
rect 113 451 129 485
rect 163 451 179 485
rect 113 417 179 451
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 113 315 129 349
rect 163 315 179 349
rect 113 265 179 315
rect 213 485 267 527
rect 213 451 223 485
rect 257 451 267 485
rect 213 417 267 451
rect 213 383 223 417
rect 257 383 267 417
rect 213 349 267 383
rect 213 315 223 349
rect 257 315 267 349
rect 213 299 267 315
rect 301 485 367 492
rect 301 451 317 485
rect 351 451 367 485
rect 301 417 367 451
rect 301 383 317 417
rect 351 383 367 417
rect 301 349 367 383
rect 401 485 455 527
rect 401 451 411 485
rect 445 451 455 485
rect 401 417 455 451
rect 401 383 411 417
rect 445 383 455 417
rect 401 367 455 383
rect 489 485 555 492
rect 489 451 505 485
rect 539 451 555 485
rect 489 417 555 451
rect 489 383 505 417
rect 539 383 555 417
rect 301 315 317 349
rect 351 333 367 349
rect 489 349 555 383
rect 589 485 643 527
rect 589 451 599 485
rect 633 451 643 485
rect 589 417 643 451
rect 589 383 599 417
rect 633 383 643 417
rect 589 367 643 383
rect 677 485 743 492
rect 677 451 693 485
rect 727 451 743 485
rect 677 417 743 451
rect 677 383 693 417
rect 727 383 743 417
rect 489 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 677 349 743 383
rect 777 485 831 527
rect 777 451 787 485
rect 821 451 831 485
rect 777 417 831 451
rect 777 383 787 417
rect 821 383 831 417
rect 777 367 831 383
rect 677 333 693 349
rect 539 315 693 333
rect 727 333 743 349
rect 727 315 815 333
rect 301 299 815 315
rect 17 249 79 265
rect 17 215 37 249
rect 71 215 79 249
rect 17 143 79 215
rect 113 249 678 265
rect 113 215 288 249
rect 322 215 356 249
rect 390 215 424 249
rect 458 215 492 249
rect 526 215 560 249
rect 594 215 628 249
rect 662 215 678 249
rect 29 93 79 109
rect 29 59 35 93
rect 69 59 79 93
rect 29 17 79 59
rect 113 106 179 215
rect 749 181 815 299
rect 301 147 815 181
rect 113 72 129 106
rect 163 72 179 106
rect 113 53 179 72
rect 213 106 267 122
rect 213 72 223 106
rect 257 72 267 106
rect 213 17 267 72
rect 301 106 367 147
rect 301 72 317 106
rect 351 72 367 106
rect 301 51 367 72
rect 401 97 455 113
rect 401 63 411 97
rect 445 63 455 97
rect 401 17 455 63
rect 489 106 555 147
rect 489 72 505 106
rect 539 72 555 106
rect 489 51 555 72
rect 589 97 643 113
rect 589 63 599 97
rect 633 63 643 97
rect 589 17 643 63
rect 677 106 743 147
rect 677 72 693 106
rect 727 72 743 106
rect 677 51 743 72
rect 777 97 831 113
rect 777 63 787 97
rect 821 63 831 97
rect 777 17 831 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel corelocali s 29 153 63 187 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel corelocali s 765 221 799 255 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel corelocali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel nbase s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 clkbuf_6
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3353952
string GDS_START 3346728
<< end >>
