magic
tech sky130A
magscale 1 2
timestamp 1601050075
<< locali >>
rect 25 224 110 426
rect 493 364 559 547
rect 493 226 551 364
rect 485 154 551 226
rect 585 162 651 310
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 22 460 72 649
rect 112 460 178 596
rect 144 330 178 460
rect 223 398 280 596
rect 316 432 363 649
rect 403 581 649 615
rect 403 398 459 581
rect 223 364 459 398
rect 593 364 649 581
rect 144 264 232 330
rect 144 162 178 264
rect 26 17 76 162
rect 112 70 178 162
rect 227 196 449 230
rect 227 70 277 196
rect 313 17 379 158
rect 415 120 449 196
rect 415 70 640 120
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel locali s 585 162 651 310 6 A
port 1 nsew signal input
rlabel locali s 25 224 110 426 6 TE_B
port 2 nsew signal input
rlabel locali s 493 364 559 547 6 Z
port 3 nsew signal output
rlabel locali s 493 226 551 364 6 Z
port 3 nsew signal output
rlabel locali s 485 154 551 226 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -49 672 49 8 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 617 672 715 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 2349900
string GDS_START 2342954
<< end >>
