magic
tech sky130A
magscale 1 2
timestamp 1599588232
<< locali >>
rect 123 368 277 430
rect 17 334 277 368
rect 17 200 51 334
rect 313 330 359 430
rect 491 342 843 376
rect 491 330 525 342
rect 313 300 415 330
rect 85 264 415 300
rect 457 264 525 330
rect 85 234 140 264
rect 619 236 743 308
rect 310 200 576 230
rect 17 196 576 200
rect 17 166 376 196
rect 21 66 87 132
rect 310 70 376 166
rect 510 70 576 196
rect 777 56 843 342
<< obsli1 >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 498 73 600
rect 113 532 367 596
rect 407 498 457 596
rect 23 464 457 498
rect 495 512 561 600
rect 595 546 661 649
rect 701 512 751 600
rect 495 478 751 512
rect 23 402 89 464
rect 407 444 457 464
rect 788 444 841 596
rect 407 410 841 444
rect 407 364 457 410
rect 121 17 276 120
rect 410 17 476 162
rect 610 17 676 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< obsli1c >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 616 50 617
rect 0 49 50 50
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel locali s 619 236 743 308 6 A
port 1 nsew signal input
rlabel locali s 777 56 843 342 6 B
port 2 nsew signal input
rlabel locali s 491 342 843 376 6 B
port 2 nsew signal input
rlabel locali s 491 330 525 342 6 B
port 2 nsew signal input
rlabel locali s 457 264 525 330 6 B
port 2 nsew signal input
rlabel locali s 313 330 359 430 6 C
port 3 nsew signal input
rlabel locali s 313 300 415 330 6 C
port 3 nsew signal input
rlabel locali s 85 264 415 300 6 C
port 3 nsew signal input
rlabel locali s 85 234 140 264 6 C
port 3 nsew signal input
rlabel locali s 21 66 87 132 6 D
port 4 nsew signal input
rlabel locali s 510 70 576 196 6 Y
port 5 nsew signal output
rlabel locali s 310 200 576 230 6 Y
port 5 nsew signal output
rlabel locali s 310 70 376 166 6 Y
port 5 nsew signal output
rlabel locali s 123 368 277 430 6 Y
port 5 nsew signal output
rlabel locali s 17 334 277 368 6 Y
port 5 nsew signal output
rlabel locali s 17 200 51 334 6 Y
port 5 nsew signal output
rlabel locali s 17 196 576 200 6 Y
port 5 nsew signal output
rlabel locali s 17 166 376 196 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -49 864 49 8 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 50 50 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 616 50 666 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 617 864 715 6 VPWR
port 9 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE /pdks/sky130A/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string GDS_END 1677912
string GDS_START 1669792
<< end >>
