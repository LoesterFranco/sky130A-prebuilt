magic
tech sky130A
magscale 1 2
timestamp 1604502723
<< locali >>
rect 121 257 187 341
rect 85 215 187 257
rect 231 289 485 341
rect 231 182 341 289
rect 231 145 475 182
rect 231 51 297 145
rect 409 51 475 145
rect 836 215 1064 255
rect 1108 215 1271 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 409 87 493
rect 127 443 203 527
rect 315 443 391 527
rect 503 443 579 527
rect 17 375 563 409
rect 17 291 87 375
rect 17 171 51 291
rect 529 323 563 375
rect 623 393 657 493
rect 710 427 760 527
rect 807 459 1053 493
rect 807 427 865 459
rect 917 393 966 425
rect 623 359 966 393
rect 529 289 641 323
rect 375 216 563 250
rect 17 53 109 171
rect 153 17 187 181
rect 341 17 375 111
rect 529 179 563 216
rect 597 249 641 289
rect 597 215 687 249
rect 749 179 787 359
rect 917 289 966 359
rect 1019 333 1053 459
rect 1087 367 1163 527
rect 1207 333 1262 493
rect 1019 291 1262 333
rect 529 129 787 179
rect 831 145 1262 181
rect 831 95 881 145
rect 513 17 579 95
rect 621 51 881 95
rect 925 17 959 111
rect 993 51 1069 145
rect 1113 17 1147 111
rect 1181 53 1262 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 1108 215 1271 255 6 A1
port 1 nsew signal input
rlabel locali s 836 215 1064 255 6 A2
port 2 nsew signal input
rlabel locali s 121 257 187 341 6 B1_N
port 3 nsew signal input
rlabel locali s 85 215 187 257 6 B1_N
port 3 nsew signal input
rlabel locali s 409 51 475 145 6 X
port 4 nsew signal output
rlabel locali s 231 289 485 341 6 X
port 4 nsew signal output
rlabel locali s 231 182 341 289 6 X
port 4 nsew signal output
rlabel locali s 231 145 475 182 6 X
port 4 nsew signal output
rlabel locali s 231 51 297 145 6 X
port 4 nsew signal output
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 6 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string LEFview TRUE
string GDS_FILE /home/aag/sky130A-prebuilt/sky130A/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 1070004
string GDS_START 1060508
<< end >>
